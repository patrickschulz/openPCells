.SUBCKT DFFNQR CLK D Q RST VDD VSS
*.PININFO CLK:I D:I RST:I Q:O VDD:B VSS:B
MN53 net9 RST VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN63 mq_x VSS mq_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN46 Q qx VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 analog=0 
+ acv_opt=-1.0
MN45 net4 qx qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN52 net7 RST VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN32 net6 clkb VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN65 qf_x VSS qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN59 qx VSS VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN22 net5 clkbb VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN23 net5 clkb net5 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN24 mq D net5 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN26 clkbb VSS VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN39 mq_x clkb qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN25 clkb VSS VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN60 mq VSS mq VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM9 clkb CLK VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN44 qx qf_x net9 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM11 mq_x mq net7 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN42 net4 clkbb VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM8 net6 clkbb net6 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MMMMMMM6 net6 mq_x mq VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN43 net4 clkb net4 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN64 qf_x clkbb qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM10 clkbb clkb VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MP63 VDD VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP61 mq_x VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP13 mq D net2 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP12 net2 clkb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP11 VDD clkbb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP53 mq_x RST VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP46 qx qf_x VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP64 mq VDD mq VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP47 Q qx VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 analog=0 
+ acv_opt=-1.0
MP54 qx RST VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP33 VDD clkb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP45 qf_x qx net3 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP44 VDD clkbb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP40 mq_x clkbb qf_x VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM31 mq_x mq VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM27 mq mq_x net29 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MMMMMMM26 VDD clkbb net29 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MP65 mq_x clkb mq_x VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP43 VDD clkb net3 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM30 clkbb clkb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MMMMMMM29 clkb CLK VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP66 qf_x VDD qf_x VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP14 clkb VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP20 clkbb VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
.ENDS

