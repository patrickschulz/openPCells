* Created by KLayout

* cell register
* pin SUBSTRATE
.SUBCKT register 2
* net 2 SUBSTRATE
* device instance $1 r0 *1 44.25,1.2 slvtpfet
M$1 1 107 67 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $2 r0 *1 44.75,1.2 slvtpfet
M$2 67 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $3 r0 *1 45.25,1.2 slvtpfet
M$3 1 67 54 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $4 r0 *1 45.75,1.2 slvtpfet
M$4 54 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $5 r0 *1 46.25,1.2 slvtpfet
M$5 1 67 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $6 r0 *1 46.75,1.2 slvtpfet
M$6 1 54 24 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $7 r0 *1 47.25,1.2 slvtpfet
M$7 24 107 57 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $8 r0 *1 47.75,1.2 slvtpfet
M$8 57 1 57 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $9 r0 *1 48.25,1.2 slvtpfet
M$9 57 91 25 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $10 r0 *1 48.75,1.2 slvtpfet
M$10 25 67 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $11 r0 *1 49.25,1.2 slvtpfet
M$11 1 54 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $12 r0 *1 49.75,1.2 slvtpfet
M$12 1 57 91 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $13 r0 *1 50.25,1.2 slvtpfet
M$13 91 54 91 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $14 r0 *1 50.75,1.2 slvtpfet
M$14 91 67 59 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $15 r0 *1 51.25,1.2 slvtpfet
M$15 59 1 59 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $16 r0 *1 51.75,1.2 slvtpfet
M$16 59 92 21 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $17 r0 *1 52.25,1.2 slvtpfet
M$17 21 54 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $19 r0 *1 53.25,1.2 slvtpfet
M$19 1 59 92 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $20 r0 *1 53.75,1.2 slvtpfet
M$20 92 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $21 r0 *1 54.25,1.2 slvtpfet
M$21 1 92 106 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $22 r0 *1 54.75,1.2 slvtpfet
M$22 106 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $23 r0 *1 55.25,1.2 slvtpfet
M$23 1 106 44 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $24 r0 *1 55.75,1.2 slvtpfet
M$24 44 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $25 r0 *1 56.25,1.2 slvtpfet
M$25 1 44 45 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $26 r0 *1 56.75,1.2 slvtpfet
M$26 45 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $27 r0 *1 57.25,1.2 slvtpfet
M$27 1 44 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $28 r0 *1 57.75,1.2 slvtpfet
M$28 1 45 20 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $29 r0 *1 58.25,1.2 slvtpfet
M$29 20 106 47 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $30 r0 *1 58.75,1.2 slvtpfet
M$30 47 1 47 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $31 r0 *1 59.25,1.2 slvtpfet
M$31 47 88 19 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $32 r0 *1 59.75,1.2 slvtpfet
M$32 19 44 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $33 r0 *1 60.25,1.2 slvtpfet
M$33 1 45 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $34 r0 *1 60.75,1.2 slvtpfet
M$34 1 47 88 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $35 r0 *1 61.25,1.2 slvtpfet
M$35 88 45 88 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $36 r0 *1 61.75,1.2 slvtpfet
M$36 88 44 50 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $37 r0 *1 62.25,1.2 slvtpfet
M$37 50 1 50 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $38 r0 *1 62.75,1.2 slvtpfet
M$38 50 89 18 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $39 r0 *1 63.25,1.2 slvtpfet
M$39 18 45 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $41 r0 *1 64.25,1.2 slvtpfet
M$41 1 50 89 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $42 r0 *1 64.75,1.2 slvtpfet
M$42 89 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $43 r0 *1 65.25,1.2 slvtpfet
M$43 1 89 105 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $44 r0 *1 65.75,1.2 slvtpfet
M$44 105 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $45 r0 *1 66.25,1.2 slvtpfet
M$45 1 105 68 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $46 r0 *1 66.75,1.2 slvtpfet
M$46 68 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $47 r0 *1 67.25,1.2 slvtpfet
M$47 1 68 40 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $48 r0 *1 67.75,1.2 slvtpfet
M$48 40 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $49 r0 *1 68.25,1.2 slvtpfet
M$49 1 68 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $50 r0 *1 68.75,1.2 slvtpfet
M$50 1 40 5 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $51 r0 *1 69.25,1.2 slvtpfet
M$51 5 105 42 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $52 r0 *1 69.75,1.2 slvtpfet
M$52 42 1 42 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $53 r0 *1 70.25,1.2 slvtpfet
M$53 42 83 4 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $54 r0 *1 70.75,1.2 slvtpfet
M$54 4 68 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $55 r0 *1 71.25,1.2 slvtpfet
M$55 1 40 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $56 r0 *1 71.75,1.2 slvtpfet
M$56 1 42 83 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $57 r0 *1 72.25,1.2 slvtpfet
M$57 83 40 83 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $58 r0 *1 72.75,1.2 slvtpfet
M$58 83 68 28 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $59 r0 *1 73.25,1.2 slvtpfet
M$59 28 1 28 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $60 r0 *1 73.75,1.2 slvtpfet
M$60 28 84 3 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $61 r0 *1 74.25,1.2 slvtpfet
M$61 3 40 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $63 r0 *1 75.25,1.2 slvtpfet
M$63 1 28 84 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $64 r0 *1 75.75,1.2 slvtpfet
M$64 84 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $65 r0 *1 76.25,1.2 slvtpfet
M$65 1 84 104 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $66 r0 *1 76.75,1.2 slvtpfet
M$66 104 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $67 r0 *1 77.25,1.2 slvtpfet
M$67 1 104 30 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $68 r0 *1 77.75,1.2 slvtpfet
M$68 30 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $69 r0 *1 78.25,1.2 slvtpfet
M$69 1 30 31 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $70 r0 *1 78.75,1.2 slvtpfet
M$70 31 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $71 r0 *1 79.25,1.2 slvtpfet
M$71 1 30 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $72 r0 *1 79.75,1.2 slvtpfet
M$72 1 31 8 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $73 r0 *1 80.25,1.2 slvtpfet
M$73 8 104 33 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $74 r0 *1 80.75,1.2 slvtpfet
M$74 33 1 33 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $75 r0 *1 81.25,1.2 slvtpfet
M$75 33 85 7 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $76 r0 *1 81.75,1.2 slvtpfet
M$76 7 30 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $77 r0 *1 82.25,1.2 slvtpfet
M$77 1 31 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $78 r0 *1 82.75,1.2 slvtpfet
M$78 1 33 85 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $79 r0 *1 83.25,1.2 slvtpfet
M$79 85 31 85 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $80 r0 *1 83.75,1.2 slvtpfet
M$80 85 30 52 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $81 r0 *1 84.25,1.2 slvtpfet
M$81 52 1 52 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $82 r0 *1 84.75,1.2 slvtpfet
M$82 52 90 6 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $83 r0 *1 85.25,1.2 slvtpfet
M$83 6 31 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $85 r0 *1 86.25,1.2 slvtpfet
M$85 1 52 90 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $86 r0 *1 86.75,1.2 slvtpfet
M$86 90 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $87 r0 *1 87.25,1.2 slvtpfet
M$87 1 90 56 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $88 r0 *1 87.75,1.2 slvtpfet
M$88 56 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U PD=2.8U
* device instance $89 r0 *1 0.25,1.2 slvtpfet
M$89 1 102 100 101 slvtpfet L=0.2U W=1U AS=0.4P AD=0.15P PS=2.8U PD=1.3U
* device instance $90 r0 *1 0.75,1.2 slvtpfet
M$90 100 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $91 r0 *1 1.25,1.2 slvtpfet
M$91 1 100 80 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $92 r0 *1 1.75,1.2 slvtpfet
M$92 80 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $93 r0 *1 2.25,1.2 slvtpfet
M$93 1 100 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $94 r0 *1 2.75,1.2 slvtpfet
M$94 1 80 14 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $95 r0 *1 3.25,1.2 slvtpfet
M$95 14 99 78 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $96 r0 *1 3.75,1.2 slvtpfet
M$96 78 1 78 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $97 r0 *1 4.25,1.2 slvtpfet
M$97 78 98 10 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $98 r0 *1 4.75,1.2 slvtpfet
M$98 10 100 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $99 r0 *1 5.25,1.2 slvtpfet
M$99 1 80 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $100 r0 *1 5.75,1.2 slvtpfet
M$100 1 78 98 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $101 r0 *1 6.25,1.2 slvtpfet
M$101 98 80 98 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $102 r0 *1 6.75,1.2 slvtpfet
M$102 98 100 66 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $103 r0 *1 7.25,1.2 slvtpfet
M$103 66 1 66 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $104 r0 *1 7.75,1.2 slvtpfet
M$104 66 93 9 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $105 r0 *1 8.25,1.2 slvtpfet
M$105 9 80 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $107 r0 *1 9.25,1.2 slvtpfet
M$107 1 66 93 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $108 r0 *1 9.75,1.2 slvtpfet
M$108 93 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $109 r0 *1 10.25,1.2 slvtpfet
M$109 1 93 103 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $110 r0 *1 10.75,1.2 slvtpfet
M$110 103 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $111 r0 *1 11.25,1.2 slvtpfet
M$111 1 103 64 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $112 r0 *1 11.75,1.2 slvtpfet
M$112 64 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $113 r0 *1 12.25,1.2 slvtpfet
M$113 1 64 63 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $114 r0 *1 12.75,1.2 slvtpfet
M$114 63 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $115 r0 *1 13.25,1.2 slvtpfet
M$115 1 64 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $116 r0 *1 13.75,1.2 slvtpfet
M$116 1 63 17 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $117 r0 *1 14.25,1.2 slvtpfet
M$117 17 103 61 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $118 r0 *1 14.75,1.2 slvtpfet
M$118 61 1 61 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $119 r0 *1 15.25,1.2 slvtpfet
M$119 61 95 16 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $120 r0 *1 15.75,1.2 slvtpfet
M$120 16 64 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $121 r0 *1 16.25,1.2 slvtpfet
M$121 1 63 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $122 r0 *1 16.75,1.2 slvtpfet
M$122 1 61 95 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $123 r0 *1 17.25,1.2 slvtpfet
M$123 95 63 95 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $124 r0 *1 17.75,1.2 slvtpfet
M$124 95 64 70 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $125 r0 *1 18.25,1.2 slvtpfet
M$125 70 1 70 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $126 r0 *1 18.75,1.2 slvtpfet
M$126 70 94 15 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $127 r0 *1 19.25,1.2 slvtpfet
M$127 15 63 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $129 r0 *1 20.25,1.2 slvtpfet
M$129 1 70 94 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $130 r0 *1 20.75,1.2 slvtpfet
M$130 94 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $131 r0 *1 21.25,1.2 slvtpfet
M$131 1 94 109 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $132 r0 *1 21.75,1.2 slvtpfet
M$132 109 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $133 r0 *1 22.25,1.2 slvtpfet
M$133 1 109 48 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $134 r0 *1 22.75,1.2 slvtpfet
M$134 48 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $135 r0 *1 23.25,1.2 slvtpfet
M$135 1 48 39 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $136 r0 *1 23.75,1.2 slvtpfet
M$136 39 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $137 r0 *1 24.25,1.2 slvtpfet
M$137 1 48 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $138 r0 *1 24.75,1.2 slvtpfet
M$138 1 39 26 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $139 r0 *1 25.25,1.2 slvtpfet
M$139 26 109 37 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $140 r0 *1 25.75,1.2 slvtpfet
M$140 37 1 37 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $141 r0 *1 26.25,1.2 slvtpfet
M$141 37 87 23 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $142 r0 *1 26.75,1.2 slvtpfet
M$142 23 48 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $143 r0 *1 27.25,1.2 slvtpfet
M$143 1 39 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $144 r0 *1 27.75,1.2 slvtpfet
M$144 1 37 87 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $145 r0 *1 28.25,1.2 slvtpfet
M$145 87 39 87 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $146 r0 *1 28.75,1.2 slvtpfet
M$146 87 48 36 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $147 r0 *1 29.25,1.2 slvtpfet
M$147 36 1 36 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $148 r0 *1 29.75,1.2 slvtpfet
M$148 36 86 22 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $149 r0 *1 30.25,1.2 slvtpfet
M$149 22 39 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $151 r0 *1 31.25,1.2 slvtpfet
M$151 1 36 86 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $152 r0 *1 31.75,1.2 slvtpfet
M$152 86 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $153 r0 *1 32.25,1.2 slvtpfet
M$153 1 86 108 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $154 r0 *1 32.75,1.2 slvtpfet
M$154 108 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $155 r0 *1 33.25,1.2 slvtpfet
M$155 1 108 81 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $156 r0 *1 33.75,1.2 slvtpfet
M$156 81 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $157 r0 *1 34.25,1.2 slvtpfet
M$157 1 81 82 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $158 r0 *1 34.75,1.2 slvtpfet
M$158 82 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $159 r0 *1 35.25,1.2 slvtpfet
M$159 1 81 1 101 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $160 r0 *1 35.75,1.2 slvtpfet
M$160 1 82 13 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $161 r0 *1 36.25,1.2 slvtpfet
M$161 13 108 75 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $162 r0 *1 36.75,1.2 slvtpfet
M$162 75 1 75 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $163 r0 *1 37.25,1.2 slvtpfet
M$163 75 97 12 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $164 r0 *1 37.75,1.2 slvtpfet
M$164 12 81 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $165 r0 *1 38.25,1.2 slvtpfet
M$165 1 82 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $166 r0 *1 38.75,1.2 slvtpfet
M$166 1 75 97 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $167 r0 *1 39.25,1.2 slvtpfet
M$167 97 82 97 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $168 r0 *1 39.75,1.2 slvtpfet
M$168 97 81 73 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $169 r0 *1 40.25,1.2 slvtpfet
M$169 73 1 73 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $170 r0 *1 40.75,1.2 slvtpfet
M$170 73 96 11 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $171 r0 *1 41.25,1.2 slvtpfet
M$171 11 82 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $173 r0 *1 42.25,1.2 slvtpfet
M$173 1 73 96 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $174 r0 *1 42.75,1.2 slvtpfet
M$174 96 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $175 r0 *1 43.25,1.2 slvtpfet
M$175 1 96 107 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $176 r0 *1 43.75,1.2 slvtpfet
M$176 107 1 1 101 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $177 r0 *1 44.25,-1.2 slvtnfet
M$177 1 107 67 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $178 r0 *1 44.75,-1.2 slvtnfet
M$178 67 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $179 r0 *1 45.25,-1.2 slvtnfet
M$179 1 67 54 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $180 r0 *1 45.75,-1.2 slvtnfet
M$180 54 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $181 r0 *1 46.25,-1.2 slvtnfet
M$181 1 67 53 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $182 r0 *1 46.75,-1.2 slvtnfet
M$182 53 54 53 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $183 r0 *1 47.25,-1.2 slvtnfet
M$183 53 107 57 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $184 r0 *1 47.75,-1.2 slvtnfet
M$184 57 1 57 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $185 r0 *1 48.25,-1.2 slvtnfet
M$185 57 91 58 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $186 r0 *1 48.75,-1.2 slvtnfet
M$186 58 67 58 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $187 r0 *1 49.25,-1.2 slvtnfet
M$187 58 54 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $188 r0 *1 49.75,-1.2 slvtnfet
M$188 1 57 91 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $189 r0 *1 50.25,-1.2 slvtnfet
M$189 91 54 59 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $190 r0 *1 50.75,-1.2 slvtnfet
M$190 59 67 59 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $191 r0 *1 51.25,-1.2 slvtnfet
M$191 59 1 59 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $192 r0 *1 51.75,-1.2 slvtnfet
M$192 59 92 60 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $193 r0 *1 52.25,-1.2 slvtnfet
M$193 60 54 60 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $194 r0 *1 52.75,-1.2 slvtnfet
M$194 60 67 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $195 r0 *1 53.25,-1.2 slvtnfet
M$195 1 59 92 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $196 r0 *1 53.75,-1.2 slvtnfet
M$196 92 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $197 r0 *1 54.25,-1.2 slvtnfet
M$197 1 92 106 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $198 r0 *1 54.75,-1.2 slvtnfet
M$198 106 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $199 r0 *1 55.25,-1.2 slvtnfet
M$199 1 106 44 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $200 r0 *1 55.75,-1.2 slvtnfet
M$200 44 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $201 r0 *1 56.25,-1.2 slvtnfet
M$201 1 44 45 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $202 r0 *1 56.75,-1.2 slvtnfet
M$202 45 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $203 r0 *1 57.25,-1.2 slvtnfet
M$203 1 44 46 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $204 r0 *1 57.75,-1.2 slvtnfet
M$204 46 45 46 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $205 r0 *1 58.25,-1.2 slvtnfet
M$205 46 106 47 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $206 r0 *1 58.75,-1.2 slvtnfet
M$206 47 1 47 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $207 r0 *1 59.25,-1.2 slvtnfet
M$207 47 88 49 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $208 r0 *1 59.75,-1.2 slvtnfet
M$208 49 44 49 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $209 r0 *1 60.25,-1.2 slvtnfet
M$209 49 45 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $210 r0 *1 60.75,-1.2 slvtnfet
M$210 1 47 88 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $211 r0 *1 61.25,-1.2 slvtnfet
M$211 88 45 50 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $212 r0 *1 61.75,-1.2 slvtnfet
M$212 50 44 50 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $213 r0 *1 62.25,-1.2 slvtnfet
M$213 50 1 50 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $214 r0 *1 62.75,-1.2 slvtnfet
M$214 50 89 51 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $215 r0 *1 63.25,-1.2 slvtnfet
M$215 51 45 51 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $216 r0 *1 63.75,-1.2 slvtnfet
M$216 51 44 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $217 r0 *1 64.25,-1.2 slvtnfet
M$217 1 50 89 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $218 r0 *1 64.75,-1.2 slvtnfet
M$218 89 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $219 r0 *1 65.25,-1.2 slvtnfet
M$219 1 89 105 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $220 r0 *1 65.75,-1.2 slvtnfet
M$220 105 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $221 r0 *1 66.25,-1.2 slvtnfet
M$221 1 105 68 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $222 r0 *1 66.75,-1.2 slvtnfet
M$222 68 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $223 r0 *1 67.25,-1.2 slvtnfet
M$223 1 68 40 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $224 r0 *1 67.75,-1.2 slvtnfet
M$224 40 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $225 r0 *1 68.25,-1.2 slvtnfet
M$225 1 68 41 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $226 r0 *1 68.75,-1.2 slvtnfet
M$226 41 40 41 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $227 r0 *1 69.25,-1.2 slvtnfet
M$227 41 105 42 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $228 r0 *1 69.75,-1.2 slvtnfet
M$228 42 1 42 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $229 r0 *1 70.25,-1.2 slvtnfet
M$229 42 83 27 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $230 r0 *1 70.75,-1.2 slvtnfet
M$230 27 68 27 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $231 r0 *1 71.25,-1.2 slvtnfet
M$231 27 40 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $232 r0 *1 71.75,-1.2 slvtnfet
M$232 1 42 83 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $233 r0 *1 72.25,-1.2 slvtnfet
M$233 83 40 28 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $234 r0 *1 72.75,-1.2 slvtnfet
M$234 28 68 28 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $235 r0 *1 73.25,-1.2 slvtnfet
M$235 28 1 28 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $236 r0 *1 73.75,-1.2 slvtnfet
M$236 28 84 29 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $237 r0 *1 74.25,-1.2 slvtnfet
M$237 29 40 29 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $238 r0 *1 74.75,-1.2 slvtnfet
M$238 29 68 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $239 r0 *1 75.25,-1.2 slvtnfet
M$239 1 28 84 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $240 r0 *1 75.75,-1.2 slvtnfet
M$240 84 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $241 r0 *1 76.25,-1.2 slvtnfet
M$241 1 84 104 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $242 r0 *1 76.75,-1.2 slvtnfet
M$242 104 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $243 r0 *1 77.25,-1.2 slvtnfet
M$243 1 104 30 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $244 r0 *1 77.75,-1.2 slvtnfet
M$244 30 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $245 r0 *1 78.25,-1.2 slvtnfet
M$245 1 30 31 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $246 r0 *1 78.75,-1.2 slvtnfet
M$246 31 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $247 r0 *1 79.25,-1.2 slvtnfet
M$247 1 30 32 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $248 r0 *1 79.75,-1.2 slvtnfet
M$248 32 31 32 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $249 r0 *1 80.25,-1.2 slvtnfet
M$249 32 104 33 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $250 r0 *1 80.75,-1.2 slvtnfet
M$250 33 1 33 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $251 r0 *1 81.25,-1.2 slvtnfet
M$251 33 85 34 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $252 r0 *1 81.75,-1.2 slvtnfet
M$252 34 30 34 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $253 r0 *1 82.25,-1.2 slvtnfet
M$253 34 31 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $254 r0 *1 82.75,-1.2 slvtnfet
M$254 1 33 85 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $255 r0 *1 83.25,-1.2 slvtnfet
M$255 85 31 52 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $256 r0 *1 83.75,-1.2 slvtnfet
M$256 52 30 52 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $257 r0 *1 84.25,-1.2 slvtnfet
M$257 52 1 52 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $258 r0 *1 84.75,-1.2 slvtnfet
M$258 52 90 55 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $259 r0 *1 85.25,-1.2 slvtnfet
M$259 55 31 55 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $260 r0 *1 85.75,-1.2 slvtnfet
M$260 55 30 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $261 r0 *1 86.25,-1.2 slvtnfet
M$261 1 52 90 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $262 r0 *1 86.75,-1.2 slvtnfet
M$262 90 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $263 r0 *1 87.25,-1.2 slvtnfet
M$263 1 90 56 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $264 r0 *1 87.75,-1.2 slvtnfet
M$264 56 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U PD=2.8U
* device instance $265 r0 *1 0.25,-1.2 slvtnfet
M$265 1 102 100 2 slvtnfet L=0.2U W=1U AS=0.4P AD=0.15P PS=2.8U PD=1.3U
* device instance $266 r0 *1 0.75,-1.2 slvtnfet
M$266 100 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $267 r0 *1 1.25,-1.2 slvtnfet
M$267 1 100 80 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $268 r0 *1 1.75,-1.2 slvtnfet
M$268 80 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $269 r0 *1 2.25,-1.2 slvtnfet
M$269 1 100 79 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $270 r0 *1 2.75,-1.2 slvtnfet
M$270 79 80 79 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $271 r0 *1 3.25,-1.2 slvtnfet
M$271 79 99 78 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $272 r0 *1 3.75,-1.2 slvtnfet
M$272 78 1 78 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $273 r0 *1 4.25,-1.2 slvtnfet
M$273 78 98 77 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $274 r0 *1 4.75,-1.2 slvtnfet
M$274 77 100 77 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $275 r0 *1 5.25,-1.2 slvtnfet
M$275 77 80 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $276 r0 *1 5.75,-1.2 slvtnfet
M$276 1 78 98 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $277 r0 *1 6.25,-1.2 slvtnfet
M$277 98 80 66 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $278 r0 *1 6.75,-1.2 slvtnfet
M$278 66 100 66 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $279 r0 *1 7.25,-1.2 slvtnfet
M$279 66 1 66 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $280 r0 *1 7.75,-1.2 slvtnfet
M$280 66 93 65 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $281 r0 *1 8.25,-1.2 slvtnfet
M$281 65 80 65 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $282 r0 *1 8.75,-1.2 slvtnfet
M$282 65 100 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $283 r0 *1 9.25,-1.2 slvtnfet
M$283 1 66 93 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $284 r0 *1 9.75,-1.2 slvtnfet
M$284 93 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $285 r0 *1 10.25,-1.2 slvtnfet
M$285 1 93 103 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $286 r0 *1 10.75,-1.2 slvtnfet
M$286 103 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $287 r0 *1 11.25,-1.2 slvtnfet
M$287 1 103 64 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $288 r0 *1 11.75,-1.2 slvtnfet
M$288 64 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $289 r0 *1 12.25,-1.2 slvtnfet
M$289 1 64 63 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $290 r0 *1 12.75,-1.2 slvtnfet
M$290 63 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $291 r0 *1 13.25,-1.2 slvtnfet
M$291 1 64 62 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $292 r0 *1 13.75,-1.2 slvtnfet
M$292 62 63 62 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $293 r0 *1 14.25,-1.2 slvtnfet
M$293 62 103 61 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $294 r0 *1 14.75,-1.2 slvtnfet
M$294 61 1 61 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $295 r0 *1 15.25,-1.2 slvtnfet
M$295 61 95 71 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $296 r0 *1 15.75,-1.2 slvtnfet
M$296 71 64 71 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $297 r0 *1 16.25,-1.2 slvtnfet
M$297 71 63 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $298 r0 *1 16.75,-1.2 slvtnfet
M$298 1 61 95 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $299 r0 *1 17.25,-1.2 slvtnfet
M$299 95 63 70 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $300 r0 *1 17.75,-1.2 slvtnfet
M$300 70 64 70 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $301 r0 *1 18.25,-1.2 slvtnfet
M$301 70 1 70 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $302 r0 *1 18.75,-1.2 slvtnfet
M$302 70 94 69 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $303 r0 *1 19.25,-1.2 slvtnfet
M$303 69 63 69 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $304 r0 *1 19.75,-1.2 slvtnfet
M$304 69 64 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $305 r0 *1 20.25,-1.2 slvtnfet
M$305 1 70 94 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $306 r0 *1 20.75,-1.2 slvtnfet
M$306 94 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $307 r0 *1 21.25,-1.2 slvtnfet
M$307 1 94 109 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $308 r0 *1 21.75,-1.2 slvtnfet
M$308 109 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $309 r0 *1 22.25,-1.2 slvtnfet
M$309 1 109 48 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $310 r0 *1 22.75,-1.2 slvtnfet
M$310 48 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $311 r0 *1 23.25,-1.2 slvtnfet
M$311 1 48 39 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $312 r0 *1 23.75,-1.2 slvtnfet
M$312 39 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $313 r0 *1 24.25,-1.2 slvtnfet
M$313 1 48 38 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $314 r0 *1 24.75,-1.2 slvtnfet
M$314 38 39 38 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $315 r0 *1 25.25,-1.2 slvtnfet
M$315 38 109 37 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $316 r0 *1 25.75,-1.2 slvtnfet
M$316 37 1 37 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $317 r0 *1 26.25,-1.2 slvtnfet
M$317 37 87 43 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $318 r0 *1 26.75,-1.2 slvtnfet
M$318 43 48 43 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $319 r0 *1 27.25,-1.2 slvtnfet
M$319 43 39 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $320 r0 *1 27.75,-1.2 slvtnfet
M$320 1 37 87 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $321 r0 *1 28.25,-1.2 slvtnfet
M$321 87 39 36 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $322 r0 *1 28.75,-1.2 slvtnfet
M$322 36 48 36 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $323 r0 *1 29.25,-1.2 slvtnfet
M$323 36 1 36 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $324 r0 *1 29.75,-1.2 slvtnfet
M$324 36 86 35 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $325 r0 *1 30.25,-1.2 slvtnfet
M$325 35 39 35 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $326 r0 *1 30.75,-1.2 slvtnfet
M$326 35 48 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $327 r0 *1 31.25,-1.2 slvtnfet
M$327 1 36 86 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $328 r0 *1 31.75,-1.2 slvtnfet
M$328 86 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $329 r0 *1 32.25,-1.2 slvtnfet
M$329 1 86 108 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $330 r0 *1 32.75,-1.2 slvtnfet
M$330 108 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $331 r0 *1 33.25,-1.2 slvtnfet
M$331 1 108 81 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $332 r0 *1 33.75,-1.2 slvtnfet
M$332 81 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $333 r0 *1 34.25,-1.2 slvtnfet
M$333 1 81 82 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $334 r0 *1 34.75,-1.2 slvtnfet
M$334 82 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $335 r0 *1 35.25,-1.2 slvtnfet
M$335 1 81 76 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $336 r0 *1 35.75,-1.2 slvtnfet
M$336 76 82 76 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $337 r0 *1 36.25,-1.2 slvtnfet
M$337 76 108 75 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $338 r0 *1 36.75,-1.2 slvtnfet
M$338 75 1 75 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $339 r0 *1 37.25,-1.2 slvtnfet
M$339 75 97 74 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $340 r0 *1 37.75,-1.2 slvtnfet
M$340 74 81 74 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $341 r0 *1 38.25,-1.2 slvtnfet
M$341 74 82 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $342 r0 *1 38.75,-1.2 slvtnfet
M$342 1 75 97 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $343 r0 *1 39.25,-1.2 slvtnfet
M$343 97 82 73 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $344 r0 *1 39.75,-1.2 slvtnfet
M$344 73 81 73 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $345 r0 *1 40.25,-1.2 slvtnfet
M$345 73 1 73 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $346 r0 *1 40.75,-1.2 slvtnfet
M$346 73 96 72 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $347 r0 *1 41.25,-1.2 slvtnfet
M$347 72 82 72 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $348 r0 *1 41.75,-1.2 slvtnfet
M$348 72 81 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $349 r0 *1 42.25,-1.2 slvtnfet
M$349 1 73 96 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $350 r0 *1 42.75,-1.2 slvtnfet
M$350 96 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $351 r0 *1 43.25,-1.2 slvtnfet
M$351 1 96 107 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $352 r0 *1 43.75,-1.2 slvtnfet
M$352 107 1 1 2 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
.ENDS register
