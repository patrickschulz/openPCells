* Created by KLayout

* cell nor_gate
* pin SUBSTRATE
.SUBCKT nor_gate 8
* net 8 SUBSTRATE
* device instance $1 r0 *1 -0.25,1.2 slvtpfet
M$1 2 3 7 6 slvtpfet L=0.2U W=1U AS=0.4P AD=0.15P PS=2.8U PD=1.3U
* device instance $2 r0 *1 0.25,1.2 slvtpfet
M$2 7 5 4 6 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $3 r0 *1 0.75,1.2 slvtpfet
M$3 4 2 2 6 slvtpfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U PD=2.8U
* device instance $4 r0 *1 -0.25,-1.2 slvtnfet
M$4 1 3 4 8 slvtnfet L=0.2U W=1U AS=0.4P AD=0.15P PS=2.8U PD=1.3U
* device instance $5 r0 *1 0.25,-1.2 slvtnfet
M$5 4 5 1 8 slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $6 r0 *1 0.75,-1.2 slvtnfet
M$6 1 1 1 8 slvtnfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U PD=2.8U
.ENDS nor_gate
