* Created by KLayout

* cell register
* pin SUBSTRATE
.SUBCKT register SUBSTRATE
* device instance $1 r0 *1 42.25,1.2 slvtpfet
M$1 \$1 \$1 \$I426 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $3 r0 *1 43.25,1.2 slvtpfet
M$3 \$1 \$I426 \$I463 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $4 r0 *1 43.75,1.2 slvtpfet
M$4 \$I463 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $5 r0 *1 44.25,1.2 slvtpfet
M$5 \$1 \$I426 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $6 r0 *1 44.75,1.2 slvtpfet
M$6 \$1 \$I463 \$I1110 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $7 r0 *1 45.25,1.2 slvtpfet
M$7 \$I1110 \$1 \$I454 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $8 r0 *1 45.75,1.2 slvtpfet
M$8 \$I454 \$1 \$I454 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $9 r0 *1 46.25,1.2 slvtpfet
M$9 \$I454 \$I122 \$I1107 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $10 r0 *1 46.75,1.2 slvtpfet
M$10 \$I1107 \$I426 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $11 r0 *1 47.25,1.2 slvtpfet
M$11 \$1 \$I463 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $12 r0 *1 47.75,1.2 slvtpfet
M$12 \$1 \$I454 \$I122 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $13 r0 *1 48.25,1.2 slvtpfet
M$13 \$I122 \$I463 \$I122 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $14 r0 *1 48.75,1.2 slvtpfet
M$14 \$I122 \$I426 \$I448 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $15 r0 *1 49.25,1.2 slvtpfet
M$15 \$I448 \$1 \$I448 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $16 r0 *1 49.75,1.2 slvtpfet
M$16 \$I448 \$I128 \$I1134 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $17 r0 *1 50.25,1.2 slvtpfet
M$17 \$I1134 \$I463 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $19 r0 *1 51.25,1.2 slvtpfet
M$19 \$1 \$I448 \$I128 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $20 r0 *1 51.75,1.2 slvtpfet
M$20 \$I128 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $21 r0 *1 52.25,1.2 slvtpfet
M$21 \$1 \$I128 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $22 r0 *1 52.75,1.2 slvtpfet
M$22 \$1 \$1 \$I490 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $24 r0 *1 53.75,1.2 slvtpfet
M$24 \$1 \$I490 \$I488 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $25 r0 *1 54.25,1.2 slvtpfet
M$25 \$I488 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $26 r0 *1 54.75,1.2 slvtpfet
M$26 \$1 \$I490 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $27 r0 *1 55.25,1.2 slvtpfet
M$27 \$1 \$I488 \$I1145 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $28 r0 *1 55.75,1.2 slvtpfet
M$28 \$I1145 \$1 \$I471 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $29 r0 *1 56.25,1.2 slvtpfet
M$29 \$I471 \$1 \$I471 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $30 r0 *1 56.75,1.2 slvtpfet
M$30 \$I471 \$I152 \$I1148 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $31 r0 *1 57.25,1.2 slvtpfet
M$31 \$I1148 \$I490 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $32 r0 *1 57.75,1.2 slvtpfet
M$32 \$1 \$I488 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $33 r0 *1 58.25,1.2 slvtpfet
M$33 \$1 \$I471 \$I152 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $34 r0 *1 58.75,1.2 slvtpfet
M$34 \$I152 \$I488 \$I152 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $35 r0 *1 59.25,1.2 slvtpfet
M$35 \$I152 \$I490 \$I478 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $36 r0 *1 59.75,1.2 slvtpfet
M$36 \$I478 \$1 \$I478 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $37 r0 *1 60.25,1.2 slvtpfet
M$37 \$I478 \$I145 \$I1155 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $38 r0 *1 60.75,1.2 slvtpfet
M$38 \$I1155 \$I488 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $40 r0 *1 61.75,1.2 slvtpfet
M$40 \$1 \$I478 \$I145 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $41 r0 *1 62.25,1.2 slvtpfet
M$41 \$I145 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $42 r0 *1 62.75,1.2 slvtpfet
M$42 \$1 \$I145 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $43 r0 *1 63.25,1.2 slvtpfet
M$43 \$1 \$1 \$I423 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $45 r0 *1 64.25,1.2 slvtpfet
M$45 \$1 \$I423 \$I501 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $46 r0 *1 64.75,1.2 slvtpfet
M$46 \$I501 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $47 r0 *1 65.25,1.2 slvtpfet
M$47 \$1 \$I423 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $48 r0 *1 65.75,1.2 slvtpfet
M$48 \$1 \$I501 \$I1251 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $49 r0 *1 66.25,1.2 slvtpfet
M$49 \$I1251 \$1 \$I509 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $50 r0 *1 66.75,1.2 slvtpfet
M$50 \$I509 \$1 \$I509 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $51 r0 *1 67.25,1.2 slvtpfet
M$51 \$I509 \$I215 \$I1259 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $52 r0 *1 67.75,1.2 slvtpfet
M$52 \$I1259 \$I423 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $53 r0 *1 68.25,1.2 slvtpfet
M$53 \$1 \$I501 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $54 r0 *1 68.75,1.2 slvtpfet
M$54 \$1 \$I509 \$I215 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $55 r0 *1 69.25,1.2 slvtpfet
M$55 \$I215 \$I501 \$I215 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $56 r0 *1 69.75,1.2 slvtpfet
M$56 \$I215 \$I423 \$I541 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $57 r0 *1 70.25,1.2 slvtpfet
M$57 \$I541 \$1 \$I541 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $58 r0 *1 70.75,1.2 slvtpfet
M$58 \$I541 \$I208 \$I1260 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $59 r0 *1 71.25,1.2 slvtpfet
M$59 \$I1260 \$I501 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $61 r0 *1 72.25,1.2 slvtpfet
M$61 \$1 \$I541 \$I208 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $62 r0 *1 72.75,1.2 slvtpfet
M$62 \$I208 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $63 r0 *1 73.25,1.2 slvtpfet
M$63 \$1 \$I208 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $64 r0 *1 73.75,1.2 slvtpfet
M$64 \$1 \$1 \$I532 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $66 r0 *1 74.75,1.2 slvtpfet
M$66 \$1 \$I532 \$I530 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $67 r0 *1 75.25,1.2 slvtpfet
M$67 \$I530 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $68 r0 *1 75.75,1.2 slvtpfet
M$68 \$1 \$I532 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $69 r0 *1 76.25,1.2 slvtpfet
M$69 \$1 \$I530 \$I1227 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $70 r0 *1 76.75,1.2 slvtpfet
M$70 \$I1227 \$1 \$I526 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $71 r0 *1 77.25,1.2 slvtpfet
M$71 \$I526 \$1 \$I526 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $72 r0 *1 77.75,1.2 slvtpfet
M$72 \$I526 \$I194 \$I1230 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $73 r0 *1 78.25,1.2 slvtpfet
M$73 \$I1230 \$I532 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $74 r0 *1 78.75,1.2 slvtpfet
M$74 \$1 \$I530 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $75 r0 *1 79.25,1.2 slvtpfet
M$75 \$1 \$I526 \$I194 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $76 r0 *1 79.75,1.2 slvtpfet
M$76 \$I194 \$I530 \$I194 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $77 r0 *1 80.25,1.2 slvtpfet
M$77 \$I194 \$I532 \$I467 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $78 r0 *1 80.75,1.2 slvtpfet
M$78 \$I467 \$1 \$I467 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $79 r0 *1 81.25,1.2 slvtpfet
M$79 \$I467 \$I130 \$I1237 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $80 r0 *1 81.75,1.2 slvtpfet
M$80 \$I1237 \$I530 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $82 r0 *1 82.75,1.2 slvtpfet
M$82 \$1 \$I467 \$I130 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $83 r0 *1 83.25,1.2 slvtpfet
M$83 \$I130 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $84 r0 *1 83.75,1.2 slvtpfet
M$84 \$1 \$I130 \$2 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U PD=2.8U
* device instance $85 r0 *1 0.25,1.2 slvtpfet
M$85 \$1 \$I21 \$I50 \$I35 slvtpfet L=0.2U W=1U AS=0.4P AD=0.15P PS=2.8U PD=1.3U
* device instance $86 r0 *1 0.75,1.2 slvtpfet
M$86 \$I50 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $87 r0 *1 1.25,1.2 slvtpfet
M$87 \$1 \$I50 \$I387 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $88 r0 *1 1.75,1.2 slvtpfet
M$88 \$I387 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $89 r0 *1 2.25,1.2 slvtpfet
M$89 \$1 \$I50 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $90 r0 *1 2.75,1.2 slvtpfet
M$90 \$1 \$I387 \$I1186 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $91 r0 *1 3.25,1.2 slvtpfet
M$91 \$I1186 \$I61 \$I391 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $92 r0 *1 3.75,1.2 slvtpfet
M$92 \$I391 \$1 \$I391 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $93 r0 *1 4.25,1.2 slvtpfet
M$93 \$I391 \$I51 \$I1211 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $94 r0 *1 4.75,1.2 slvtpfet
M$94 \$I1211 \$I50 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $95 r0 *1 5.25,1.2 slvtpfet
M$95 \$1 \$I387 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $96 r0 *1 5.75,1.2 slvtpfet
M$96 \$1 \$I391 \$I51 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $97 r0 *1 6.25,1.2 slvtpfet
M$97 \$I51 \$I387 \$I51 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $98 r0 *1 6.75,1.2 slvtpfet
M$98 \$I51 \$I50 \$I430 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $99 r0 *1 7.25,1.2 slvtpfet
M$99 \$I430 \$1 \$I430 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $100 r0 *1 7.75,1.2 slvtpfet
M$100 \$I430 \$I103 \$I1174 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $101 r0 *1 8.25,1.2 slvtpfet
M$101 \$I1174 \$I387 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $103 r0 *1 9.25,1.2 slvtpfet
M$103 \$1 \$I430 \$I103 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $104 r0 *1 9.75,1.2 slvtpfet
M$104 \$I103 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $105 r0 *1 10.25,1.2 slvtpfet
M$105 \$1 \$I103 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $106 r0 *1 10.75,1.2 slvtpfet
M$106 \$1 \$1 \$I439 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $108 r0 *1 11.75,1.2 slvtpfet
M$108 \$1 \$I439 \$I441 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $109 r0 *1 12.25,1.2 slvtpfet
M$109 \$I441 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $110 r0 *1 12.75,1.2 slvtpfet
M$110 \$1 \$I439 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $111 r0 *1 13.25,1.2 slvtpfet
M$111 \$1 \$I441 \$I1169 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $112 r0 *1 13.75,1.2 slvtpfet
M$112 \$I1169 \$1 \$I419 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $113 r0 *1 14.25,1.2 slvtpfet
M$113 \$I419 \$1 \$I419 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $114 r0 *1 14.75,1.2 slvtpfet
M$114 \$I419 \$I81 \$I1172 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $115 r0 *1 15.25,1.2 slvtpfet
M$115 \$I1172 \$I439 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $116 r0 *1 15.75,1.2 slvtpfet
M$116 \$1 \$I441 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $117 r0 *1 16.25,1.2 slvtpfet
M$117 \$1 \$I419 \$I81 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $118 r0 *1 16.75,1.2 slvtpfet
M$118 \$I81 \$I441 \$I81 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $119 r0 *1 17.25,1.2 slvtpfet
M$119 \$I81 \$I439 \$I415 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $120 r0 *1 17.75,1.2 slvtpfet
M$120 \$I415 \$1 \$I415 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $121 r0 *1 18.25,1.2 slvtpfet
M$121 \$I415 \$I88 \$I1179 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $122 r0 *1 18.75,1.2 slvtpfet
M$122 \$I1179 \$I441 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $124 r0 *1 19.75,1.2 slvtpfet
M$124 \$1 \$I415 \$I88 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $125 r0 *1 20.25,1.2 slvtpfet
M$125 \$I88 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $126 r0 *1 20.75,1.2 slvtpfet
M$126 \$1 \$I88 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $127 r0 *1 21.25,1.2 slvtpfet
M$127 \$1 \$1 \$I484 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $129 r0 *1 22.25,1.2 slvtpfet
M$129 \$1 \$I484 \$I504 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $130 r0 *1 22.75,1.2 slvtpfet
M$130 \$I504 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $131 r0 *1 23.25,1.2 slvtpfet
M$131 \$1 \$I484 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $132 r0 *1 23.75,1.2 slvtpfet
M$132 \$1 \$I504 \$I1097 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $133 r0 *1 24.25,1.2 slvtpfet
M$133 \$I1097 \$1 \$I508 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $134 r0 *1 24.75,1.2 slvtpfet
M$134 \$I508 \$1 \$I508 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $135 r0 *1 25.25,1.2 slvtpfet
M$135 \$I508 \$I180 \$I1115 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $136 r0 *1 25.75,1.2 slvtpfet
M$136 \$I1115 \$I484 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $137 r0 *1 26.25,1.2 slvtpfet
M$137 \$1 \$I504 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $138 r0 *1 26.75,1.2 slvtpfet
M$138 \$1 \$I508 \$I180 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $139 r0 *1 27.25,1.2 slvtpfet
M$139 \$I180 \$I504 \$I180 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $140 r0 *1 27.75,1.2 slvtpfet
M$140 \$I180 \$I484 \$I514 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $141 r0 *1 28.25,1.2 slvtpfet
M$141 \$I514 \$1 \$I514 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $142 r0 *1 28.75,1.2 slvtpfet
M$142 \$I514 \$I187 \$I1122 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $143 r0 *1 29.25,1.2 slvtpfet
M$143 \$I1122 \$I504 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $145 r0 *1 30.25,1.2 slvtpfet
M$145 \$1 \$I514 \$I187 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $146 r0 *1 30.75,1.2 slvtpfet
M$146 \$I187 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $147 r0 *1 31.25,1.2 slvtpfet
M$147 \$1 \$I187 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $148 r0 *1 31.75,1.2 slvtpfet
M$148 \$1 \$1 \$I385 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $150 r0 *1 32.75,1.2 slvtpfet
M$150 \$1 \$I385 \$I382 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $151 r0 *1 33.25,1.2 slvtpfet
M$151 \$I382 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $152 r0 *1 33.75,1.2 slvtpfet
M$152 \$1 \$I385 \$1 \$I35 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $153 r0 *1 34.25,1.2 slvtpfet
M$153 \$1 \$I382 \$I1193 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $154 r0 *1 34.75,1.2 slvtpfet
M$154 \$I1193 \$1 \$I405 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $155 r0 *1 35.25,1.2 slvtpfet
M$155 \$I405 \$1 \$I405 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $156 r0 *1 35.75,1.2 slvtpfet
M$156 \$I405 \$I73 \$I1196 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $157 r0 *1 36.25,1.2 slvtpfet
M$157 \$I1196 \$I385 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $158 r0 *1 36.75,1.2 slvtpfet
M$158 \$1 \$I382 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $159 r0 *1 37.25,1.2 slvtpfet
M$159 \$1 \$I405 \$I73 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $160 r0 *1 37.75,1.2 slvtpfet
M$160 \$I73 \$I382 \$I73 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $161 r0 *1 38.25,1.2 slvtpfet
M$161 \$I73 \$I385 \$I399 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $162 r0 *1 38.75,1.2 slvtpfet
M$162 \$I399 \$1 \$I399 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $163 r0 *1 39.25,1.2 slvtpfet
M$163 \$I399 \$I66 \$I1188 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $164 r0 *1 39.75,1.2 slvtpfet
M$164 \$I1188 \$I382 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $166 r0 *1 40.75,1.2 slvtpfet
M$166 \$1 \$I399 \$I66 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $167 r0 *1 41.25,1.2 slvtpfet
M$167 \$I66 \$1 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $168 r0 *1 41.75,1.2 slvtpfet
M$168 \$1 \$I66 \$1 \$I35 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $169 r0 *1 42.25,-1.2 slvtnfet
M$169 \$1 \$1 \$I426 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $171 r0 *1 43.25,-1.2 slvtnfet
M$171 \$1 \$I426 \$I463 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $172 r0 *1 43.75,-1.2 slvtnfet
M$172 \$I463 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $173 r0 *1 44.25,-1.2 slvtnfet
M$173 \$1 \$I426 \$I465 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $174 r0 *1 44.75,-1.2 slvtnfet
M$174 \$I465 \$I463 \$I465 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $175 r0 *1 45.25,-1.2 slvtnfet
M$175 \$I465 \$1 \$I454 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $176 r0 *1 45.75,-1.2 slvtnfet
M$176 \$I454 \$1 \$I454 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $177 r0 *1 46.25,-1.2 slvtnfet
M$177 \$I454 \$I122 \$I452 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $178 r0 *1 46.75,-1.2 slvtnfet
M$178 \$I452 \$I426 \$I452 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $179 r0 *1 47.25,-1.2 slvtnfet
M$179 \$I452 \$I463 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $180 r0 *1 47.75,-1.2 slvtnfet
M$180 \$1 \$I454 \$I122 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $181 r0 *1 48.25,-1.2 slvtnfet
M$181 \$I122 \$I463 \$I448 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $182 r0 *1 48.75,-1.2 slvtnfet
M$182 \$I448 \$I426 \$I448 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $183 r0 *1 49.25,-1.2 slvtnfet
M$183 \$I448 \$1 \$I448 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $184 r0 *1 49.75,-1.2 slvtnfet
M$184 \$I448 \$I128 \$I458 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $185 r0 *1 50.25,-1.2 slvtnfet
M$185 \$I458 \$I463 \$I458 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $186 r0 *1 50.75,-1.2 slvtnfet
M$186 \$I458 \$I426 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $187 r0 *1 51.25,-1.2 slvtnfet
M$187 \$1 \$I448 \$I128 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $188 r0 *1 51.75,-1.2 slvtnfet
M$188 \$I128 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $189 r0 *1 52.25,-1.2 slvtnfet
M$189 \$1 \$I128 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $190 r0 *1 52.75,-1.2 slvtnfet
M$190 \$1 \$1 \$I490 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $192 r0 *1 53.75,-1.2 slvtnfet
M$192 \$1 \$I490 \$I488 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $193 r0 *1 54.25,-1.2 slvtnfet
M$193 \$I488 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $194 r0 *1 54.75,-1.2 slvtnfet
M$194 \$1 \$I490 \$I486 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $195 r0 *1 55.25,-1.2 slvtnfet
M$195 \$I486 \$I488 \$I486 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $196 r0 *1 55.75,-1.2 slvtnfet
M$196 \$I486 \$1 \$I471 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $197 r0 *1 56.25,-1.2 slvtnfet
M$197 \$I471 \$1 \$I471 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $198 r0 *1 56.75,-1.2 slvtnfet
M$198 \$I471 \$I152 \$I482 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $199 r0 *1 57.25,-1.2 slvtnfet
M$199 \$I482 \$I490 \$I482 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $200 r0 *1 57.75,-1.2 slvtnfet
M$200 \$I482 \$I488 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $201 r0 *1 58.25,-1.2 slvtnfet
M$201 \$1 \$I471 \$I152 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $202 r0 *1 58.75,-1.2 slvtnfet
M$202 \$I152 \$I488 \$I478 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $203 r0 *1 59.25,-1.2 slvtnfet
M$203 \$I478 \$I490 \$I478 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $204 r0 *1 59.75,-1.2 slvtnfet
M$204 \$I478 \$1 \$I478 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $205 r0 *1 60.25,-1.2 slvtnfet
M$205 \$I478 \$I145 \$I475 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $206 r0 *1 60.75,-1.2 slvtnfet
M$206 \$I475 \$I488 \$I475 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $207 r0 *1 61.25,-1.2 slvtnfet
M$207 \$I475 \$I490 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $208 r0 *1 61.75,-1.2 slvtnfet
M$208 \$1 \$I478 \$I145 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $209 r0 *1 62.25,-1.2 slvtnfet
M$209 \$I145 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $210 r0 *1 62.75,-1.2 slvtnfet
M$210 \$1 \$I145 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $211 r0 *1 63.25,-1.2 slvtnfet
M$211 \$1 \$1 \$I423 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $213 r0 *1 64.25,-1.2 slvtnfet
M$213 \$1 \$I423 \$I501 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $214 r0 *1 64.75,-1.2 slvtnfet
M$214 \$I501 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $215 r0 *1 65.25,-1.2 slvtnfet
M$215 \$1 \$I423 \$I499 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $216 r0 *1 65.75,-1.2 slvtnfet
M$216 \$I499 \$I501 \$I499 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $217 r0 *1 66.25,-1.2 slvtnfet
M$217 \$I499 \$1 \$I509 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $218 r0 *1 66.75,-1.2 slvtnfet
M$218 \$I509 \$1 \$I509 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $219 r0 *1 67.25,-1.2 slvtnfet
M$219 \$I509 \$I215 \$I545 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $220 r0 *1 67.75,-1.2 slvtnfet
M$220 \$I545 \$I423 \$I545 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $221 r0 *1 68.25,-1.2 slvtnfet
M$221 \$I545 \$I501 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $222 r0 *1 68.75,-1.2 slvtnfet
M$222 \$1 \$I509 \$I215 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $223 r0 *1 69.25,-1.2 slvtnfet
M$223 \$I215 \$I501 \$I541 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $224 r0 *1 69.75,-1.2 slvtnfet
M$224 \$I541 \$I423 \$I541 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $225 r0 *1 70.25,-1.2 slvtnfet
M$225 \$I541 \$1 \$I541 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $226 r0 *1 70.75,-1.2 slvtnfet
M$226 \$I541 \$I208 \$I538 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $227 r0 *1 71.25,-1.2 slvtnfet
M$227 \$I538 \$I501 \$I538 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $228 r0 *1 71.75,-1.2 slvtnfet
M$228 \$I538 \$I423 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $229 r0 *1 72.25,-1.2 slvtnfet
M$229 \$1 \$I541 \$I208 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $230 r0 *1 72.75,-1.2 slvtnfet
M$230 \$I208 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $231 r0 *1 73.25,-1.2 slvtnfet
M$231 \$1 \$I208 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $232 r0 *1 73.75,-1.2 slvtnfet
M$232 \$1 \$1 \$I532 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $234 r0 *1 74.75,-1.2 slvtnfet
M$234 \$1 \$I532 \$I530 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $235 r0 *1 75.25,-1.2 slvtnfet
M$235 \$I530 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $236 r0 *1 75.75,-1.2 slvtnfet
M$236 \$1 \$I532 \$I528 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $237 r0 *1 76.25,-1.2 slvtnfet
M$237 \$I528 \$I530 \$I528 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $238 r0 *1 76.75,-1.2 slvtnfet
M$238 \$I528 \$1 \$I526 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $239 r0 *1 77.25,-1.2 slvtnfet
M$239 \$I526 \$1 \$I526 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $240 r0 *1 77.75,-1.2 slvtnfet
M$240 \$I526 \$I194 \$I524 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $241 r0 *1 78.25,-1.2 slvtnfet
M$241 \$I524 \$I532 \$I524 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $242 r0 *1 78.75,-1.2 slvtnfet
M$242 \$I524 \$I530 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $243 r0 *1 79.25,-1.2 slvtnfet
M$243 \$1 \$I526 \$I194 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $244 r0 *1 79.75,-1.2 slvtnfet
M$244 \$I194 \$I530 \$I467 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $245 r0 *1 80.25,-1.2 slvtnfet
M$245 \$I467 \$I532 \$I467 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $246 r0 *1 80.75,-1.2 slvtnfet
M$246 \$I467 \$1 \$I467 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $247 r0 *1 81.25,-1.2 slvtnfet
M$247 \$I467 \$I130 \$I460 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $248 r0 *1 81.75,-1.2 slvtnfet
M$248 \$I460 \$I530 \$I460 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $249 r0 *1 82.25,-1.2 slvtnfet
M$249 \$I460 \$I532 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $250 r0 *1 82.75,-1.2 slvtnfet
M$250 \$1 \$I467 \$I130 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $251 r0 *1 83.25,-1.2 slvtnfet
M$251 \$I130 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $252 r0 *1 83.75,-1.2 slvtnfet
M$252 \$1 \$I130 \$2 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U
+ PD=2.8U
* device instance $253 r0 *1 0.25,-1.2 slvtnfet
M$253 \$1 \$I21 \$I50 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.4P AD=0.15P PS=2.8U
+ PD=1.3U
* device instance $254 r0 *1 0.75,-1.2 slvtnfet
M$254 \$I50 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $255 r0 *1 1.25,-1.2 slvtnfet
M$255 \$1 \$I50 \$I387 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $256 r0 *1 1.75,-1.2 slvtnfet
M$256 \$I387 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $257 r0 *1 2.25,-1.2 slvtnfet
M$257 \$1 \$I50 \$I389 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $258 r0 *1 2.75,-1.2 slvtnfet
M$258 \$I389 \$I387 \$I389 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $259 r0 *1 3.25,-1.2 slvtnfet
M$259 \$I389 \$I61 \$I391 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $260 r0 *1 3.75,-1.2 slvtnfet
M$260 \$I391 \$1 \$I391 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $261 r0 *1 4.25,-1.2 slvtnfet
M$261 \$I391 \$I51 \$I381 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $262 r0 *1 4.75,-1.2 slvtnfet
M$262 \$I381 \$I50 \$I381 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $263 r0 *1 5.25,-1.2 slvtnfet
M$263 \$I381 \$I387 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $264 r0 *1 5.75,-1.2 slvtnfet
M$264 \$1 \$I391 \$I51 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $265 r0 *1 6.25,-1.2 slvtnfet
M$265 \$I51 \$I387 \$I430 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $266 r0 *1 6.75,-1.2 slvtnfet
M$266 \$I430 \$I50 \$I430 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $267 r0 *1 7.25,-1.2 slvtnfet
M$267 \$I430 \$1 \$I430 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $268 r0 *1 7.75,-1.2 slvtnfet
M$268 \$I430 \$I103 \$I433 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $269 r0 *1 8.25,-1.2 slvtnfet
M$269 \$I433 \$I387 \$I433 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $270 r0 *1 8.75,-1.2 slvtnfet
M$270 \$I433 \$I50 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $271 r0 *1 9.25,-1.2 slvtnfet
M$271 \$1 \$I430 \$I103 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $272 r0 *1 9.75,-1.2 slvtnfet
M$272 \$I103 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $273 r0 *1 10.25,-1.2 slvtnfet
M$273 \$1 \$I103 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $274 r0 *1 10.75,-1.2 slvtnfet
M$274 \$1 \$1 \$I439 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $276 r0 *1 11.75,-1.2 slvtnfet
M$276 \$1 \$I439 \$I441 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $277 r0 *1 12.25,-1.2 slvtnfet
M$277 \$I441 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $278 r0 *1 12.75,-1.2 slvtnfet
M$278 \$1 \$I439 \$I443 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $279 r0 *1 13.25,-1.2 slvtnfet
M$279 \$I443 \$I441 \$I443 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $280 r0 *1 13.75,-1.2 slvtnfet
M$280 \$I443 \$1 \$I419 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $281 r0 *1 14.25,-1.2 slvtnfet
M$281 \$I419 \$1 \$I419 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $282 r0 *1 14.75,-1.2 slvtnfet
M$282 \$I419 \$I81 \$I411 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $283 r0 *1 15.25,-1.2 slvtnfet
M$283 \$I411 \$I439 \$I411 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $284 r0 *1 15.75,-1.2 slvtnfet
M$284 \$I411 \$I441 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $285 r0 *1 16.25,-1.2 slvtnfet
M$285 \$1 \$I419 \$I81 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $286 r0 *1 16.75,-1.2 slvtnfet
M$286 \$I81 \$I441 \$I415 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $287 r0 *1 17.25,-1.2 slvtnfet
M$287 \$I415 \$I439 \$I415 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $288 r0 *1 17.75,-1.2 slvtnfet
M$288 \$I415 \$1 \$I415 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $289 r0 *1 18.25,-1.2 slvtnfet
M$289 \$I415 \$I88 \$I418 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $290 r0 *1 18.75,-1.2 slvtnfet
M$290 \$I418 \$I441 \$I418 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $291 r0 *1 19.25,-1.2 slvtnfet
M$291 \$I418 \$I439 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $292 r0 *1 19.75,-1.2 slvtnfet
M$292 \$1 \$I415 \$I88 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $293 r0 *1 20.25,-1.2 slvtnfet
M$293 \$I88 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $294 r0 *1 20.75,-1.2 slvtnfet
M$294 \$1 \$I88 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $295 r0 *1 21.25,-1.2 slvtnfet
M$295 \$1 \$1 \$I484 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $297 r0 *1 22.25,-1.2 slvtnfet
M$297 \$1 \$I484 \$I504 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $298 r0 *1 22.75,-1.2 slvtnfet
M$298 \$I504 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $299 r0 *1 23.25,-1.2 slvtnfet
M$299 \$1 \$I484 \$I506 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $300 r0 *1 23.75,-1.2 slvtnfet
M$300 \$I506 \$I504 \$I506 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $301 r0 *1 24.25,-1.2 slvtnfet
M$301 \$I506 \$1 \$I508 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $302 r0 *1 24.75,-1.2 slvtnfet
M$302 \$I508 \$1 \$I508 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $303 r0 *1 25.25,-1.2 slvtnfet
M$303 \$I508 \$I180 \$I510 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $304 r0 *1 25.75,-1.2 slvtnfet
M$304 \$I510 \$I484 \$I510 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $305 r0 *1 26.25,-1.2 slvtnfet
M$305 \$I510 \$I504 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $306 r0 *1 26.75,-1.2 slvtnfet
M$306 \$1 \$I508 \$I180 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $307 r0 *1 27.25,-1.2 slvtnfet
M$307 \$I180 \$I504 \$I514 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $308 r0 *1 27.75,-1.2 slvtnfet
M$308 \$I514 \$I484 \$I514 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $309 r0 *1 28.25,-1.2 slvtnfet
M$309 \$I514 \$1 \$I514 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $310 r0 *1 28.75,-1.2 slvtnfet
M$310 \$I514 \$I187 \$I517 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $311 r0 *1 29.25,-1.2 slvtnfet
M$311 \$I517 \$I504 \$I517 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $312 r0 *1 29.75,-1.2 slvtnfet
M$312 \$I517 \$I484 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $313 r0 *1 30.25,-1.2 slvtnfet
M$313 \$1 \$I514 \$I187 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $314 r0 *1 30.75,-1.2 slvtnfet
M$314 \$I187 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $315 r0 *1 31.25,-1.2 slvtnfet
M$315 \$1 \$I187 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $316 r0 *1 31.75,-1.2 slvtnfet
M$316 \$1 \$1 \$I385 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $318 r0 *1 32.75,-1.2 slvtnfet
M$318 \$1 \$I385 \$I382 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $319 r0 *1 33.25,-1.2 slvtnfet
M$319 \$I382 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $320 r0 *1 33.75,-1.2 slvtnfet
M$320 \$1 \$I385 \$I408 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $321 r0 *1 34.25,-1.2 slvtnfet
M$321 \$I408 \$I382 \$I408 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $322 r0 *1 34.75,-1.2 slvtnfet
M$322 \$I408 \$1 \$I405 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $323 r0 *1 35.25,-1.2 slvtnfet
M$323 \$I405 \$1 \$I405 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $324 r0 *1 35.75,-1.2 slvtnfet
M$324 \$I405 \$I73 \$I403 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $325 r0 *1 36.25,-1.2 slvtnfet
M$325 \$I403 \$I385 \$I403 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $326 r0 *1 36.75,-1.2 slvtnfet
M$326 \$I403 \$I382 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $327 r0 *1 37.25,-1.2 slvtnfet
M$327 \$1 \$I405 \$I73 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $328 r0 *1 37.75,-1.2 slvtnfet
M$328 \$I73 \$I382 \$I399 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $329 r0 *1 38.25,-1.2 slvtnfet
M$329 \$I399 \$I385 \$I399 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $330 r0 *1 38.75,-1.2 slvtnfet
M$330 \$I399 \$1 \$I399 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $331 r0 *1 39.25,-1.2 slvtnfet
M$331 \$I399 \$I66 \$I396 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $332 r0 *1 39.75,-1.2 slvtnfet
M$332 \$I396 \$I382 \$I396 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $333 r0 *1 40.25,-1.2 slvtnfet
M$333 \$I396 \$I385 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $334 r0 *1 40.75,-1.2 slvtnfet
M$334 \$1 \$I399 \$I66 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $335 r0 *1 41.25,-1.2 slvtnfet
M$335 \$I66 \$1 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $336 r0 *1 41.75,-1.2 slvtnfet
M$336 \$1 \$I66 \$1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
.ENDS register
