* Created by KLayout

* cell all_cells
* pin SUBSTRATE
.SUBCKT all_cells SUBSTRATE
* device instance $1 r0 *1 41.75,1.2 slvtpfet
M$1 \$I1 \$I359 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $2 r0 *1 42.25,1.2 slvtpfet
M$2 \$I1 \$I1 \$I580 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $4 r0 *1 43.25,1.2 slvtpfet
M$4 \$I1 \$I580 \$I677 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $5 r0 *1 43.75,1.2 slvtpfet
M$5 \$I677 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U PD=1.3U
* device instance $6 r0 *1 44.25,1.2 slvtpfet
M$6 \$I1 \$I580 \$I1 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $7 r0 *1 44.75,1.2 slvtpfet
M$7 \$I1 \$I677 \$I1301 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $8 r0 *1 45.25,1.2 slvtpfet
M$8 \$I1301 \$I1 \$I589 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $9 r0 *1 45.75,1.2 slvtpfet
M$9 \$I589 \$I1 \$I589 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $10 r0 *1 46.25,1.2 slvtpfet
M$10 \$I589 \$I303 \$I1314 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $11 r0 *1 46.75,1.2 slvtpfet
M$11 \$I1314 \$I580 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $12 r0 *1 47.25,1.2 slvtpfet
M$12 \$I1 \$I677 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $13 r0 *1 47.75,1.2 slvtpfet
M$13 \$I1 \$I589 \$I303 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $14 r0 *1 48.25,1.2 slvtpfet
M$14 \$I303 \$I677 \$I303 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $15 r0 *1 48.75,1.2 slvtpfet
M$15 \$I303 \$I580 \$I583 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $16 r0 *1 49.25,1.2 slvtpfet
M$16 \$I583 \$I1 \$I583 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $17 r0 *1 49.75,1.2 slvtpfet
M$17 \$I583 \$I328 \$I1323 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $18 r0 *1 50.25,1.2 slvtpfet
M$18 \$I1323 \$I677 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $20 r0 *1 51.25,1.2 slvtpfet
M$20 \$I1 \$I583 \$I328 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $21 r0 *1 51.75,1.2 slvtpfet
M$21 \$I328 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $22 r0 *1 52.25,1.2 slvtpfet
M$22 \$I1 \$I328 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $23 r0 *1 52.75,1.2 slvtpfet
M$23 \$I1 \$I1 \$I618 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $25 r0 *1 53.75,1.2 slvtpfet
M$25 \$I1 \$I618 \$I620 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $26 r0 *1 54.25,1.2 slvtpfet
M$26 \$I620 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $27 r0 *1 54.75,1.2 slvtpfet
M$27 \$I1 \$I618 \$I1 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $28 r0 *1 55.25,1.2 slvtpfet
M$28 \$I1 \$I620 \$I1334 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $29 r0 *1 55.75,1.2 slvtpfet
M$29 \$I1334 \$I1 \$I610 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $30 r0 *1 56.25,1.2 slvtpfet
M$30 \$I610 \$I1 \$I610 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $31 r0 *1 56.75,1.2 slvtpfet
M$31 \$I610 \$I342 \$I1337 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $32 r0 *1 57.25,1.2 slvtpfet
M$32 \$I1337 \$I618 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $33 r0 *1 57.75,1.2 slvtpfet
M$33 \$I1 \$I620 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $34 r0 *1 58.25,1.2 slvtpfet
M$34 \$I1 \$I610 \$I342 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $35 r0 *1 58.75,1.2 slvtpfet
M$35 \$I342 \$I620 \$I342 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $36 r0 *1 59.25,1.2 slvtpfet
M$36 \$I342 \$I618 \$I630 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $37 r0 *1 59.75,1.2 slvtpfet
M$37 \$I630 \$I1 \$I630 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $38 r0 *1 60.25,1.2 slvtpfet
M$38 \$I630 \$I349 \$I1294 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $39 r0 *1 60.75,1.2 slvtpfet
M$39 \$I1294 \$I620 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $41 r0 *1 61.75,1.2 slvtpfet
M$41 \$I1 \$I630 \$I349 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $42 r0 *1 62.25,1.2 slvtpfet
M$42 \$I349 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $43 r0 *1 62.75,1.2 slvtpfet
M$43 \$I1 \$I349 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $44 r0 *1 63.25,1.2 slvtpfet
M$44 \$I1 \$I1 \$I573 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $46 r0 *1 64.25,1.2 slvtpfet
M$46 \$I1 \$I573 \$I653 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $47 r0 *1 64.75,1.2 slvtpfet
M$47 \$I653 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $48 r0 *1 65.25,1.2 slvtpfet
M$48 \$I1 \$I573 \$I1 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $49 r0 *1 65.75,1.2 slvtpfet
M$49 \$I1 \$I653 \$I1404 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $50 r0 *1 66.25,1.2 slvtpfet
M$50 \$I1404 \$I1 \$I680 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $51 r0 *1 66.75,1.2 slvtpfet
M$51 \$I680 \$I1 \$I680 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $52 r0 *1 67.25,1.2 slvtpfet
M$52 \$I680 \$I397 \$I1389 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $53 r0 *1 67.75,1.2 slvtpfet
M$53 \$I1389 \$I573 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $54 r0 *1 68.25,1.2 slvtpfet
M$54 \$I1 \$I653 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $55 r0 *1 68.75,1.2 slvtpfet
M$55 \$I1 \$I680 \$I397 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $56 r0 *1 69.25,1.2 slvtpfet
M$56 \$I397 \$I653 \$I397 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $57 r0 *1 69.75,1.2 slvtpfet
M$57 \$I397 \$I573 \$I674 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $58 r0 *1 70.25,1.2 slvtpfet
M$58 \$I674 \$I1 \$I674 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $59 r0 *1 70.75,1.2 slvtpfet
M$59 \$I674 \$I387 \$I1414 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $60 r0 *1 71.25,1.2 slvtpfet
M$60 \$I1414 \$I653 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $62 r0 *1 72.25,1.2 slvtpfet
M$62 \$I1 \$I674 \$I387 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $63 r0 *1 72.75,1.2 slvtpfet
M$63 \$I387 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $64 r0 *1 73.25,1.2 slvtpfet
M$64 \$I1 \$I387 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $65 r0 *1 73.75,1.2 slvtpfet
M$65 \$I1 \$I1 \$I651 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $67 r0 *1 74.75,1.2 slvtpfet
M$67 \$I1 \$I651 \$I609 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $68 r0 *1 75.25,1.2 slvtpfet
M$68 \$I609 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $69 r0 *1 75.75,1.2 slvtpfet
M$69 \$I1 \$I651 \$I1 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $70 r0 *1 76.25,1.2 slvtpfet
M$70 \$I1 \$I609 \$I1425 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $71 r0 *1 76.75,1.2 slvtpfet
M$71 \$I1425 \$I1 \$I605 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $72 r0 *1 77.25,1.2 slvtpfet
M$72 \$I605 \$I1 \$I605 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $73 r0 *1 77.75,1.2 slvtpfet
M$73 \$I605 \$I319 \$I1428 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $74 r0 *1 78.25,1.2 slvtpfet
M$74 \$I1428 \$I651 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $75 r0 *1 78.75,1.2 slvtpfet
M$75 \$I1 \$I609 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $76 r0 *1 79.25,1.2 slvtpfet
M$76 \$I1 \$I605 \$I319 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $77 r0 *1 79.75,1.2 slvtpfet
M$77 \$I319 \$I609 \$I319 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $78 r0 *1 80.25,1.2 slvtpfet
M$78 \$I319 \$I651 \$I599 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $79 r0 *1 80.75,1.2 slvtpfet
M$79 \$I599 \$I1 \$I599 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $80 r0 *1 81.25,1.2 slvtpfet
M$80 \$I599 \$I298 \$I1391 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $81 r0 *1 81.75,1.2 slvtpfet
M$81 \$I1391 \$I609 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $83 r0 *1 82.75,1.2 slvtpfet
M$83 \$I1 \$I599 \$I298 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $84 r0 *1 83.25,1.2 slvtpfet
M$84 \$I298 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $85 r0 *1 83.75,1.2 slvtpfet
M$85 \$I1 \$I298 \$I684 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.4P PS=1.3U
+ PD=2.8U
* device instance $86 r0 *1 30.25,1.2 slvtpfet
M$86 \$I1 \$I548 \$I270 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $87 r0 *1 30.75,1.2 slvtpfet
M$87 \$I270 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $88 r0 *1 31.25,1.2 slvtpfet
M$88 \$I1 \$I270 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $89 r0 *1 31.75,1.2 slvtpfet
M$89 \$I1 \$I1 \$I659 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $91 r0 *1 32.75,1.2 slvtpfet
M$91 \$I1 \$I659 \$I661 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $92 r0 *1 33.25,1.2 slvtpfet
M$92 \$I661 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $93 r0 *1 33.75,1.2 slvtpfet
M$93 \$I1 \$I659 \$I1 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $94 r0 *1 34.25,1.2 slvtpfet
M$94 \$I1 \$I661 \$I1313 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $95 r0 *1 34.75,1.2 slvtpfet
M$95 \$I1313 \$I1 \$I652 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $96 r0 *1 35.25,1.2 slvtpfet
M$96 \$I652 \$I1 \$I652 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $97 r0 *1 35.75,1.2 slvtpfet
M$97 \$I652 \$I366 \$I1365 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $98 r0 *1 36.25,1.2 slvtpfet
M$98 \$I1365 \$I659 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $99 r0 *1 36.75,1.2 slvtpfet
M$99 \$I1 \$I661 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $100 r0 *1 37.25,1.2 slvtpfet
M$100 \$I1 \$I652 \$I366 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $101 r0 *1 37.75,1.2 slvtpfet
M$101 \$I366 \$I661 \$I366 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $102 r0 *1 38.25,1.2 slvtpfet
M$102 \$I366 \$I659 \$I646 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $103 r0 *1 38.75,1.2 slvtpfet
M$103 \$I646 \$I1 \$I646 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $104 r0 *1 39.25,1.2 slvtpfet
M$104 \$I646 \$I359 \$I1372 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $105 r0 *1 39.75,1.2 slvtpfet
M$105 \$I1372 \$I661 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $107 r0 *1 40.75,1.2 slvtpfet
M$107 \$I1 \$I646 \$I359 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $108 r0 *1 41.25,1.2 slvtpfet
M$108 \$I359 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $109 r0 *1 20.75,1.2 slvtpfet
M$109 \$I1 \$I283 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $110 r0 *1 21.25,1.2 slvtpfet
M$110 \$I1 \$I1 \$I561 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $112 r0 *1 22.25,1.2 slvtpfet
M$112 \$I1 \$I561 \$I559 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $113 r0 *1 22.75,1.2 slvtpfet
M$113 \$I559 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $114 r0 *1 23.25,1.2 slvtpfet
M$114 \$I1 \$I561 \$I1 \$I4 slvtpfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U PD=2.6U
* device instance $115 r0 *1 23.75,1.2 slvtpfet
M$115 \$I1 \$I559 \$I1383 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $116 r0 *1 24.25,1.2 slvtpfet
M$116 \$I1383 \$I1 \$I552 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $117 r0 *1 24.75,1.2 slvtpfet
M$117 \$I552 \$I1 \$I552 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $118 r0 *1 25.25,1.2 slvtpfet
M$118 \$I552 \$I258 \$I1386 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $119 r0 *1 25.75,1.2 slvtpfet
M$119 \$I1386 \$I561 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $120 r0 *1 26.25,1.2 slvtpfet
M$120 \$I1 \$I559 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $121 r0 *1 26.75,1.2 slvtpfet
M$121 \$I1 \$I552 \$I258 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $122 r0 *1 27.25,1.2 slvtpfet
M$122 \$I258 \$I559 \$I258 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $123 r0 *1 27.75,1.2 slvtpfet
M$123 \$I258 \$I561 \$I548 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $124 r0 *1 28.25,1.2 slvtpfet
M$124 \$I548 \$I1 \$I548 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $125 r0 *1 28.75,1.2 slvtpfet
M$125 \$I548 \$I270 \$I1344 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $126 r0 *1 29.25,1.2 slvtpfet
M$126 \$I1344 \$I559 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $128 r0 *1 4.5,1.2 slvtpfet
M$128 \$I48 \$I1 \$I49 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $129 r0 *1 4.75,1.2 slvtpfet
M$129 \$I49 \$I1 \$I46 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $130 r0 *1 5,1.2 slvtpfet
M$130 \$I46 \$I1 \$I69 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $131 r0 *1 5.25,1.2 slvtpfet
M$131 \$I69 \$I1 \$I73 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $132 r0 *1 5.5,1.2 slvtpfet
M$132 \$I73 \$I1 \$I71 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $133 r0 *1 5.75,1.2 slvtpfet
M$133 \$I71 \$I1 \$I76 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $134 r0 *1 6,1.2 slvtpfet
M$134 \$I76 \$I1 \$I74 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $135 r0 *1 6.25,1.2 slvtpfet
M$135 \$I74 \$I1 \$I77 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $136 r0 *1 6.5,1.2 slvtpfet
M$136 \$I77 \$I1 \$I79 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $137 r0 *1 6.75,1.2 slvtpfet
M$137 \$I79 \$I1 \$I78 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $138 r0 *1 7,1.2 slvtpfet
M$138 \$I78 \$I1 \$I81 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $139 r0 *1 7.25,1.2 slvtpfet
M$139 \$I81 \$I1 \$I83 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $140 r0 *1 7.5,1.2 slvtpfet
M$140 \$I83 \$I1 \$I82 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $141 r0 *1 7.75,1.2 slvtpfet
M$141 \$I82 \$I1 \$I85 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $142 r0 *1 8,1.2 slvtpfet
M$142 \$I85 \$I1 \$I99 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $143 r0 *1 8.25,1.2 slvtpfet
M$143 \$I99 \$I1 \$I100 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $144 r0 *1 8.5,1.2 slvtpfet
M$144 \$I100 \$I1 \$I103 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $145 r0 *1 8.75,1.2 slvtpfet
M$145 \$I103 \$I1 \$I106 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $146 r0 *1 9,1.2 slvtpfet
M$146 \$I106 \$I1 \$I104 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $147 r0 *1 9.25,1.2 slvtpfet
M$147 \$I104 \$I1 \$I107 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $148 r0 *1 9.5,1.2 slvtpfet
M$148 \$I107 \$I1 \$I108 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $149 r0 *1 9.75,1.2 slvtpfet
M$149 \$I108 \$I1 \$I109 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $150 r0 *1 10,1.2 slvtpfet
M$150 \$I109 \$I1 \$I111 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $151 r0 *1 10.25,1.2 slvtpfet
M$151 \$I111 \$I1 \$I112 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $152 r0 *1 10.5,1.2 slvtpfet
M$152 \$I112 \$I1 \$I121 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $153 r0 *1 10.75,1.2 slvtpfet
M$153 \$I121 \$I1 \$I116 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $154 r0 *1 11,1.2 slvtpfet
M$154 \$I116 \$I1 \$I115 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $155 r0 *1 11.25,1.2 slvtpfet
M$155 \$I115 \$I1 \$I114 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $156 r0 *1 11.5,1.2 slvtpfet
M$156 \$I114 \$I1 \$I113 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $157 r0 *1 11.75,1.2 slvtpfet
M$157 \$I113 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.15P PS=1.05U
+ PD=1.3U
* device instance $158 r0 *1 12.25,1.2 slvtpfet
M$158 \$I1 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=4U AS=0.6P AD=0.6P PS=5.2U PD=5.2U
* device instance $160 r0 *1 13.25,1.2 slvtpfet
M$160 \$I1 \$I1 \$I1349 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $161 r0 *1 13.75,1.2 slvtpfet
M$161 \$I1349 \$I1 \$I576 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $162 r0 *1 14.25,1.2 slvtpfet
M$162 \$I576 \$I1 \$I576 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $163 r0 *1 14.75,1.2 slvtpfet
M$163 \$I576 \$I290 \$I1340 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $164 r0 *1 15.25,1.2 slvtpfet
M$164 \$I1340 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $166 r0 *1 16.25,1.2 slvtpfet
M$166 \$I1 \$I576 \$I290 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $167 r0 *1 16.75,1.2 slvtpfet
M$167 \$I290 \$I1 \$I290 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $168 r0 *1 17.25,1.2 slvtpfet
M$168 \$I290 \$I1 \$I570 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $169 r0 *1 17.75,1.2 slvtpfet
M$169 \$I570 \$I1 \$I570 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $170 r0 *1 18.25,1.2 slvtpfet
M$170 \$I570 \$I283 \$I1359 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $171 r0 *1 18.75,1.2 slvtpfet
M$171 \$I1359 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $173 r0 *1 19.75,1.2 slvtpfet
M$173 \$I1 \$I570 \$I283 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $174 r0 *1 20.25,1.2 slvtpfet
M$174 \$I283 \$I1 \$I1 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $175 r0 *1 0,1.2 slvtpfet
M$175 \$I1 \$I1 \$I6 \$I4 slvtpfet L=0.2U W=1U AS=0.15P AD=0.025P PS=1.3U
+ PD=1.05U
* device instance $176 r0 *1 0.25,1.2 slvtpfet
M$176 \$I6 \$I1 \$I7 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $177 r0 *1 0.5,1.2 slvtpfet
M$177 \$I7 \$I1 \$I20 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $178 r0 *1 0.75,1.2 slvtpfet
M$178 \$I20 \$I1 \$I21 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $179 r0 *1 1,1.2 slvtpfet
M$179 \$I21 \$I1 \$I23 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $180 r0 *1 1.25,1.2 slvtpfet
M$180 \$I23 \$I1 \$I25 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $181 r0 *1 1.5,1.2 slvtpfet
M$181 \$I25 \$I1 \$I24 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $182 r0 *1 1.75,1.2 slvtpfet
M$182 \$I24 \$I1 \$I28 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $183 r0 *1 2,1.2 slvtpfet
M$183 \$I28 \$I1 \$I26 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $184 r0 *1 2.25,1.2 slvtpfet
M$184 \$I26 \$I1 \$I29 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $185 r0 *1 2.5,1.2 slvtpfet
M$185 \$I29 \$I1 \$I30 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $186 r0 *1 2.75,1.2 slvtpfet
M$186 \$I30 \$I1 \$I31 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $187 r0 *1 3,1.2 slvtpfet
M$187 \$I31 \$I1 \$I42 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $188 r0 *1 3.25,1.2 slvtpfet
M$188 \$I42 \$I1 \$I43 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $189 r0 *1 3.5,1.2 slvtpfet
M$189 \$I43 \$I1 \$I45 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $190 r0 *1 3.75,1.2 slvtpfet
M$190 \$I45 \$I1 \$I47 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $191 r0 *1 4,1.2 slvtpfet
M$191 \$I47 \$I1 \$I44 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $192 r0 *1 4.25,1.2 slvtpfet
M$192 \$I44 \$I1 \$I48 \$I4 slvtpfet L=0.2U W=1U AS=0.025P AD=0.025P PS=1.05U
+ PD=1.05U
* device instance $193 r0 *1 41.75,-1.2 slvtnfet
M$193 \$I1 \$I359 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $194 r0 *1 42.25,-1.2 slvtnfet
M$194 \$I1 \$I1 \$I580 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $196 r0 *1 43.25,-1.2 slvtnfet
M$196 \$I1 \$I580 \$I677 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $197 r0 *1 43.75,-1.2 slvtnfet
M$197 \$I677 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $198 r0 *1 44.25,-1.2 slvtnfet
M$198 \$I1 \$I580 \$I591 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $199 r0 *1 44.75,-1.2 slvtnfet
M$199 \$I591 \$I677 \$I591 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $200 r0 *1 45.25,-1.2 slvtnfet
M$200 \$I591 \$I1 \$I589 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $201 r0 *1 45.75,-1.2 slvtnfet
M$201 \$I589 \$I1 \$I589 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $202 r0 *1 46.25,-1.2 slvtnfet
M$202 \$I589 \$I303 \$I587 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $203 r0 *1 46.75,-1.2 slvtnfet
M$203 \$I587 \$I580 \$I587 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $204 r0 *1 47.25,-1.2 slvtnfet
M$204 \$I587 \$I677 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $205 r0 *1 47.75,-1.2 slvtnfet
M$205 \$I1 \$I589 \$I303 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $206 r0 *1 48.25,-1.2 slvtnfet
M$206 \$I303 \$I677 \$I583 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $207 r0 *1 48.75,-1.2 slvtnfet
M$207 \$I583 \$I580 \$I583 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $208 r0 *1 49.25,-1.2 slvtnfet
M$208 \$I583 \$I1 \$I583 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $209 r0 *1 49.75,-1.2 slvtnfet
M$209 \$I583 \$I328 \$I612 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $210 r0 *1 50.25,-1.2 slvtnfet
M$210 \$I612 \$I677 \$I612 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $211 r0 *1 50.75,-1.2 slvtnfet
M$211 \$I612 \$I580 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $212 r0 *1 51.25,-1.2 slvtnfet
M$212 \$I1 \$I583 \$I328 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $213 r0 *1 51.75,-1.2 slvtnfet
M$213 \$I328 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $214 r0 *1 52.25,-1.2 slvtnfet
M$214 \$I1 \$I328 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $215 r0 *1 52.75,-1.2 slvtnfet
M$215 \$I1 \$I1 \$I618 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $217 r0 *1 53.75,-1.2 slvtnfet
M$217 \$I1 \$I618 \$I620 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $218 r0 *1 54.25,-1.2 slvtnfet
M$218 \$I620 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $219 r0 *1 54.75,-1.2 slvtnfet
M$219 \$I1 \$I618 \$I622 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $220 r0 *1 55.25,-1.2 slvtnfet
M$220 \$I622 \$I620 \$I622 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $221 r0 *1 55.75,-1.2 slvtnfet
M$221 \$I622 \$I1 \$I610 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $222 r0 *1 56.25,-1.2 slvtnfet
M$222 \$I610 \$I1 \$I610 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $223 r0 *1 56.75,-1.2 slvtnfet
M$223 \$I610 \$I342 \$I626 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $224 r0 *1 57.25,-1.2 slvtnfet
M$224 \$I626 \$I618 \$I626 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $225 r0 *1 57.75,-1.2 slvtnfet
M$225 \$I626 \$I620 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $226 r0 *1 58.25,-1.2 slvtnfet
M$226 \$I1 \$I610 \$I342 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $227 r0 *1 58.75,-1.2 slvtnfet
M$227 \$I342 \$I620 \$I630 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $228 r0 *1 59.25,-1.2 slvtnfet
M$228 \$I630 \$I618 \$I630 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $229 r0 *1 59.75,-1.2 slvtnfet
M$229 \$I630 \$I1 \$I630 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $230 r0 *1 60.25,-1.2 slvtnfet
M$230 \$I630 \$I349 \$I633 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $231 r0 *1 60.75,-1.2 slvtnfet
M$231 \$I633 \$I620 \$I633 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $232 r0 *1 61.25,-1.2 slvtnfet
M$232 \$I633 \$I618 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $233 r0 *1 61.75,-1.2 slvtnfet
M$233 \$I1 \$I630 \$I349 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $234 r0 *1 62.25,-1.2 slvtnfet
M$234 \$I349 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $235 r0 *1 62.75,-1.2 slvtnfet
M$235 \$I1 \$I349 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $236 r0 *1 63.25,-1.2 slvtnfet
M$236 \$I1 \$I1 \$I573 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $238 r0 *1 64.25,-1.2 slvtnfet
M$238 \$I1 \$I573 \$I653 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $239 r0 *1 64.75,-1.2 slvtnfet
M$239 \$I653 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $240 r0 *1 65.25,-1.2 slvtnfet
M$240 \$I1 \$I573 \$I639 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $241 r0 *1 65.75,-1.2 slvtnfet
M$241 \$I639 \$I653 \$I639 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $242 r0 *1 66.25,-1.2 slvtnfet
M$242 \$I639 \$I1 \$I680 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $243 r0 *1 66.75,-1.2 slvtnfet
M$243 \$I680 \$I1 \$I680 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $244 r0 *1 67.25,-1.2 slvtnfet
M$244 \$I680 \$I397 \$I681 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $245 r0 *1 67.75,-1.2 slvtnfet
M$245 \$I681 \$I573 \$I681 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $246 r0 *1 68.25,-1.2 slvtnfet
M$246 \$I681 \$I653 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $247 r0 *1 68.75,-1.2 slvtnfet
M$247 \$I1 \$I680 \$I397 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $248 r0 *1 69.25,-1.2 slvtnfet
M$248 \$I397 \$I653 \$I674 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $249 r0 *1 69.75,-1.2 slvtnfet
M$249 \$I674 \$I573 \$I674 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $250 r0 *1 70.25,-1.2 slvtnfet
M$250 \$I674 \$I1 \$I674 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $251 r0 *1 70.75,-1.2 slvtnfet
M$251 \$I674 \$I387 \$I671 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $252 r0 *1 71.25,-1.2 slvtnfet
M$252 \$I671 \$I653 \$I671 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $253 r0 *1 71.75,-1.2 slvtnfet
M$253 \$I671 \$I573 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $254 r0 *1 72.25,-1.2 slvtnfet
M$254 \$I1 \$I674 \$I387 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $255 r0 *1 72.75,-1.2 slvtnfet
M$255 \$I387 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $256 r0 *1 73.25,-1.2 slvtnfet
M$256 \$I1 \$I387 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $257 r0 *1 73.75,-1.2 slvtnfet
M$257 \$I1 \$I1 \$I651 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $259 r0 *1 74.75,-1.2 slvtnfet
M$259 \$I1 \$I651 \$I609 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $260 r0 *1 75.25,-1.2 slvtnfet
M$260 \$I609 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $261 r0 *1 75.75,-1.2 slvtnfet
M$261 \$I1 \$I651 \$I607 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $262 r0 *1 76.25,-1.2 slvtnfet
M$262 \$I607 \$I609 \$I607 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $263 r0 *1 76.75,-1.2 slvtnfet
M$263 \$I607 \$I1 \$I605 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $264 r0 *1 77.25,-1.2 slvtnfet
M$264 \$I605 \$I1 \$I605 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $265 r0 *1 77.75,-1.2 slvtnfet
M$265 \$I605 \$I319 \$I603 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $266 r0 *1 78.25,-1.2 slvtnfet
M$266 \$I603 \$I651 \$I603 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $267 r0 *1 78.75,-1.2 slvtnfet
M$267 \$I603 \$I609 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $268 r0 *1 79.25,-1.2 slvtnfet
M$268 \$I1 \$I605 \$I319 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $269 r0 *1 79.75,-1.2 slvtnfet
M$269 \$I319 \$I609 \$I599 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $270 r0 *1 80.25,-1.2 slvtnfet
M$270 \$I599 \$I651 \$I599 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $271 r0 *1 80.75,-1.2 slvtnfet
M$271 \$I599 \$I1 \$I599 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $272 r0 *1 81.25,-1.2 slvtnfet
M$272 \$I599 \$I298 \$I582 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $273 r0 *1 81.75,-1.2 slvtnfet
M$273 \$I582 \$I609 \$I582 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $274 r0 *1 82.25,-1.2 slvtnfet
M$274 \$I582 \$I651 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $275 r0 *1 82.75,-1.2 slvtnfet
M$275 \$I1 \$I599 \$I298 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $276 r0 *1 83.25,-1.2 slvtnfet
M$276 \$I298 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $277 r0 *1 83.75,-1.2 slvtnfet
M$277 \$I1 \$I298 \$I684 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.4P
+ PS=1.3U PD=2.8U
* device instance $278 r0 *1 30.25,-1.2 slvtnfet
M$278 \$I1 \$I548 \$I270 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $279 r0 *1 30.75,-1.2 slvtnfet
M$279 \$I270 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $280 r0 *1 31.25,-1.2 slvtnfet
M$280 \$I1 \$I270 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $281 r0 *1 31.75,-1.2 slvtnfet
M$281 \$I1 \$I1 \$I659 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $283 r0 *1 32.75,-1.2 slvtnfet
M$283 \$I1 \$I659 \$I661 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $284 r0 *1 33.25,-1.2 slvtnfet
M$284 \$I661 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $285 r0 *1 33.75,-1.2 slvtnfet
M$285 \$I1 \$I659 \$I663 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $286 r0 *1 34.25,-1.2 slvtnfet
M$286 \$I663 \$I661 \$I663 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $287 r0 *1 34.75,-1.2 slvtnfet
M$287 \$I663 \$I1 \$I652 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $288 r0 *1 35.25,-1.2 slvtnfet
M$288 \$I652 \$I1 \$I652 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $289 r0 *1 35.75,-1.2 slvtnfet
M$289 \$I652 \$I366 \$I650 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $290 r0 *1 36.25,-1.2 slvtnfet
M$290 \$I650 \$I659 \$I650 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $291 r0 *1 36.75,-1.2 slvtnfet
M$291 \$I650 \$I661 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $292 r0 *1 37.25,-1.2 slvtnfet
M$292 \$I1 \$I652 \$I366 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $293 r0 *1 37.75,-1.2 slvtnfet
M$293 \$I366 \$I661 \$I646 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $294 r0 *1 38.25,-1.2 slvtnfet
M$294 \$I646 \$I659 \$I646 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $295 r0 *1 38.75,-1.2 slvtnfet
M$295 \$I646 \$I1 \$I646 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $296 r0 *1 39.25,-1.2 slvtnfet
M$296 \$I646 \$I359 \$I643 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $297 r0 *1 39.75,-1.2 slvtnfet
M$297 \$I643 \$I661 \$I643 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $298 r0 *1 40.25,-1.2 slvtnfet
M$298 \$I643 \$I659 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $299 r0 *1 40.75,-1.2 slvtnfet
M$299 \$I1 \$I646 \$I359 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $300 r0 *1 41.25,-1.2 slvtnfet
M$300 \$I359 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $301 r0 *1 20.75,-1.2 slvtnfet
M$301 \$I1 \$I283 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $302 r0 *1 21.25,-1.2 slvtnfet
M$302 \$I1 \$I1 \$I561 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $304 r0 *1 22.25,-1.2 slvtnfet
M$304 \$I1 \$I561 \$I559 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $305 r0 *1 22.75,-1.2 slvtnfet
M$305 \$I559 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $306 r0 *1 23.25,-1.2 slvtnfet
M$306 \$I1 \$I561 \$I556 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $307 r0 *1 23.75,-1.2 slvtnfet
M$307 \$I556 \$I559 \$I556 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $308 r0 *1 24.25,-1.2 slvtnfet
M$308 \$I556 \$I1 \$I552 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $309 r0 *1 24.75,-1.2 slvtnfet
M$309 \$I552 \$I1 \$I552 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $310 r0 *1 25.25,-1.2 slvtnfet
M$310 \$I552 \$I258 \$I542 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $311 r0 *1 25.75,-1.2 slvtnfet
M$311 \$I542 \$I561 \$I542 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $312 r0 *1 26.25,-1.2 slvtnfet
M$312 \$I542 \$I559 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $313 r0 *1 26.75,-1.2 slvtnfet
M$313 \$I1 \$I552 \$I258 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $314 r0 *1 27.25,-1.2 slvtnfet
M$314 \$I258 \$I559 \$I548 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $315 r0 *1 27.75,-1.2 slvtnfet
M$315 \$I548 \$I561 \$I548 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $316 r0 *1 28.25,-1.2 slvtnfet
M$316 \$I548 \$I1 \$I548 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $317 r0 *1 28.75,-1.2 slvtnfet
M$317 \$I548 \$I270 \$I554 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $318 r0 *1 29.25,-1.2 slvtnfet
M$318 \$I554 \$I559 \$I554 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $319 r0 *1 29.75,-1.2 slvtnfet
M$319 \$I554 \$I561 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $320 r0 *1 4.5,-1.2 slvtnfet
M$320 \$I39 \$I1 \$I41 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $321 r0 *1 4.75,-1.2 slvtnfet
M$321 \$I41 \$I1 \$I40 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $322 r0 *1 5,-1.2 slvtnfet
M$322 \$I40 \$I1 \$I57 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $323 r0 *1 5.25,-1.2 slvtnfet
M$323 \$I57 \$I1 \$I59 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $324 r0 *1 5.5,-1.2 slvtnfet
M$324 \$I59 \$I1 \$I58 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $325 r0 *1 5.75,-1.2 slvtnfet
M$325 \$I58 \$I1 \$I61 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $326 r0 *1 6,-1.2 slvtnfet
M$326 \$I61 \$I1 \$I60 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $327 r0 *1 6.25,-1.2 slvtnfet
M$327 \$I60 \$I1 \$I64 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $328 r0 *1 6.5,-1.2 slvtnfet
M$328 \$I64 \$I1 \$I63 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $329 r0 *1 6.75,-1.2 slvtnfet
M$329 \$I63 \$I1 \$I67 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $330 r0 *1 7,-1.2 slvtnfet
M$330 \$I67 \$I1 \$I66 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $331 r0 *1 7.25,-1.2 slvtnfet
M$331 \$I66 \$I1 \$I68 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $332 r0 *1 7.5,-1.2 slvtnfet
M$332 \$I68 \$I1 \$I65 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $333 r0 *1 7.75,-1.2 slvtnfet
M$333 \$I65 \$I1 \$I62 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $334 r0 *1 8,-1.2 slvtnfet
M$334 \$I62 \$I1 \$I97 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $335 r0 *1 8.25,-1.2 slvtnfet
M$335 \$I97 \$I1 \$I98 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $336 r0 *1 8.5,-1.2 slvtnfet
M$336 \$I98 \$I1 \$I96 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $337 r0 *1 8.75,-1.2 slvtnfet
M$337 \$I96 \$I1 \$I94 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $338 r0 *1 9,-1.2 slvtnfet
M$338 \$I94 \$I1 \$I95 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $339 r0 *1 9.25,-1.2 slvtnfet
M$339 \$I95 \$I1 \$I93 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $340 r0 *1 9.5,-1.2 slvtnfet
M$340 \$I93 \$I1 \$I92 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $341 r0 *1 9.75,-1.2 slvtnfet
M$341 \$I92 \$I1 \$I91 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $342 r0 *1 10,-1.2 slvtnfet
M$342 \$I91 \$I1 \$I90 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $343 r0 *1 10.25,-1.2 slvtnfet
M$343 \$I90 \$I1 \$I89 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $344 r0 *1 10.5,-1.2 slvtnfet
M$344 \$I89 \$I1 \$I122 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $345 r0 *1 10.75,-1.2 slvtnfet
M$345 \$I122 \$I1 \$I120 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $346 r0 *1 11,-1.2 slvtnfet
M$346 \$I120 \$I1 \$I119 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $347 r0 *1 11.25,-1.2 slvtnfet
M$347 \$I119 \$I1 \$I118 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $348 r0 *1 11.5,-1.2 slvtnfet
M$348 \$I118 \$I1 \$I117 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $349 r0 *1 11.75,-1.2 slvtnfet
M$349 \$I117 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.15P
+ PS=1.05U PD=1.3U
* device instance $350 r0 *1 12.25,-1.2 slvtnfet
M$350 \$I1 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $351 r0 *1 12.75,-1.2 slvtnfet
M$351 \$I1 \$I1 \$I578 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $352 r0 *1 13.25,-1.2 slvtnfet
M$352 \$I578 \$I1 \$I578 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $353 r0 *1 13.75,-1.2 slvtnfet
M$353 \$I578 \$I1 \$I576 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $354 r0 *1 14.25,-1.2 slvtnfet
M$354 \$I576 \$I1 \$I576 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $355 r0 *1 14.75,-1.2 slvtnfet
M$355 \$I576 \$I290 \$I574 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $356 r0 *1 15.25,-1.2 slvtnfet
M$356 \$I574 \$I1 \$I574 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $357 r0 *1 15.75,-1.2 slvtnfet
M$357 \$I574 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $358 r0 *1 16.25,-1.2 slvtnfet
M$358 \$I1 \$I576 \$I290 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $359 r0 *1 16.75,-1.2 slvtnfet
M$359 \$I290 \$I1 \$I570 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $360 r0 *1 17.25,-1.2 slvtnfet
M$360 \$I570 \$I1 \$I570 SUBSTRATE slvtnfet L=0.2U W=2U AS=0.3P AD=0.3P PS=2.6U
+ PD=2.6U
* device instance $362 r0 *1 18.25,-1.2 slvtnfet
M$362 \$I570 \$I283 \$I567 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $363 r0 *1 18.75,-1.2 slvtnfet
M$363 \$I567 \$I1 \$I567 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $364 r0 *1 19.25,-1.2 slvtnfet
M$364 \$I567 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $365 r0 *1 19.75,-1.2 slvtnfet
M$365 \$I1 \$I570 \$I283 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P
+ PS=1.3U PD=1.3U
* device instance $366 r0 *1 20.25,-1.2 slvtnfet
M$366 \$I283 \$I1 \$I1 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.15P PS=1.3U
+ PD=1.3U
* device instance $367 r0 *1 0,-1.2 slvtnfet
M$367 \$I1 \$I1 \$I2 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.15P AD=0.025P PS=1.3U
+ PD=1.05U
* device instance $368 r0 *1 0.25,-1.2 slvtnfet
M$368 \$I2 \$I1 \$I3 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $369 r0 *1 0.5,-1.2 slvtnfet
M$369 \$I3 \$I1 \$I16 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $370 r0 *1 0.75,-1.2 slvtnfet
M$370 \$I16 \$I1 \$I15 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $371 r0 *1 1,-1.2 slvtnfet
M$371 \$I15 \$I1 \$I17 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $372 r0 *1 1.25,-1.2 slvtnfet
M$372 \$I17 \$I1 \$I18 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $373 r0 *1 1.5,-1.2 slvtnfet
M$373 \$I18 \$I1 \$I19 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $374 r0 *1 1.75,-1.2 slvtnfet
M$374 \$I19 \$I1 \$I13 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $375 r0 *1 2,-1.2 slvtnfet
M$375 \$I13 \$I1 \$I14 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $376 r0 *1 2.25,-1.2 slvtnfet
M$376 \$I14 \$I1 \$I12 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $377 r0 *1 2.5,-1.2 slvtnfet
M$377 \$I12 \$I1 \$I11 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $378 r0 *1 2.75,-1.2 slvtnfet
M$378 \$I11 \$I1 \$I10 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $379 r0 *1 3,-1.2 slvtnfet
M$379 \$I10 \$I1 \$I34 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $380 r0 *1 3.25,-1.2 slvtnfet
M$380 \$I34 \$I1 \$I35 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $381 r0 *1 3.5,-1.2 slvtnfet
M$381 \$I35 \$I1 \$I37 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $382 r0 *1 3.75,-1.2 slvtnfet
M$382 \$I37 \$I1 \$I38 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $383 r0 *1 4,-1.2 slvtnfet
M$383 \$I38 \$I1 \$I36 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
* device instance $384 r0 *1 4.25,-1.2 slvtnfet
M$384 \$I36 \$I1 \$I39 SUBSTRATE slvtnfet L=0.2U W=1U AS=0.025P AD=0.025P
+ PS=1.05U PD=1.05U
.ENDS all_cells
