.SUBCKT DFFNQS CLK D Q SET VDD VSS
*.PININFO CLK:I D:I SET:I Q:O VDD:B VSS:B
MN51 net1 VSS net1 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN50 net0 VSS net0 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN49 net1 SET VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN46 Q qx VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 analog=0 
+ acv_opt=-1.0
MN47 qx VSS VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN45 net4 qx qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN48 net0 SET VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN32 net6 clkb net0 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN41 qf_x VSS qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN22 net5 clkbb VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN23 net5 clkb net5 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN24 mq D net5 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN26 clkbb VSS VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN39 mq_x clkb qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN25 clkb VSS VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN28 mq VSS mq VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN40 qf_x clkbb qf_x VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM9 clkb CLK VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN44 qx qf_x VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM11 mq_x mq VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN42 net4 clkbb net1 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM8 net6 clkbb net6 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MMMMMMM6 net6 mq_x mq VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MN43 net4 clkb net4 VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM10 clkbb clkb VSS VSS slvtnfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MP52 qf_x VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP51 mq VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP13 mq D net2 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP12 net2 clkb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP11 VDD clkbb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP48 qx VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP46 qx qf_x VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP47 Q qx VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 analog=0 
+ acv_opt=-1.0
MP49 mq SET VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP50 qf_x SET VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP33 VDD clkb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP42 qf_x VDD qf_x VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP45 qf_x qx net3 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP44 VDD clkbb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP40 mq_x clkbb qf_x VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM31 mq_x mq VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM27 mq mq_x net29 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MMMMMMM26 VDD clkbb net29 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MP43 VDD clkb net3 VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MMMMMMM30 clkbb clkb VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 
+ ngcon=1 analog=0 acv_opt=-1.0
MMMMMMM29 clkb CLK VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP22 mq VDD mq VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP14 clkb VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP41 mq_x clkb mq_x VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
MP20 clkbb VDD VDD VSS slvtpfet m=1 w=300n l=40n nf=1 p_la=0 ulp=0 ngcon=1 
+ analog=0 acv_opt=-1.0
.ENDS

